
        // PE 0, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[0][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[0][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[0][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[0][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[0][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[0][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[0][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[0][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[0][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[0][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[0][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[0][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[0][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[0][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[0][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[0][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[0][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[0][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[0][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[0][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[0][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[0][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[0][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[0][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[0][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[0][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[0][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[0][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[0][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[0][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[0][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[0][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[0][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[0][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[0][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[0][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[0][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[0][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[0][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[0][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[0][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[0][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[0][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[0][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[0][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[0][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[0][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[0][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[0][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[0][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[0][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[0][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[0][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[0][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[0][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[0][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[0][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[0][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[0][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[0][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[0][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[0][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[0][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[0][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[0][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[0][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[0][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[0][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[0][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[0][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[0][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[0][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[0][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[0][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[0][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[0][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[0][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[0][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[0][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[0][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[0][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[0][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[0][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[0][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[0][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[0][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[0][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[0][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[0][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[0][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[0][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[0][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[0][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[0][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[0][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[0][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[0][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[0][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[0][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[0][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[0][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[0][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[0][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[0][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[0][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[0][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[0][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[0][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[0][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[0][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[0][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[0][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[0][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[0][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[0][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[0][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[0][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[0][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[0][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[0][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[0][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[0][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[0][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[0][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[0][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[0][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[0][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[0][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[0][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[0][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[0][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[0][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[0][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[0][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[0][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[0][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[0][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[0][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[0][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[0][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[0][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[0][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[0][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[0][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[0][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[0][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[0][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[0][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[0][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[0][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[0][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[0][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[0][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[0][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[0][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[0][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[0][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[0][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[0][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[0][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[0][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[0][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[0][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[0][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[0][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[0][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[0][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[0][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[0][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[0][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[0][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[0][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[0][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[0][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[0][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[0][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[0][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[0][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[0][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[0][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[0][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[0][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[0][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[0][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[0][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[0][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 0, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[0][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[0][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[0][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[0][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[0][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[0].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[0][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[1][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[1][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[1][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[1][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[1][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[1][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[1][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[1][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[1][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[1][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[1][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[1][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[1][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[1][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[1][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[1][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[1][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[1][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[1][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[1][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[1][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[1][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[1][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[1][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[1][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[1][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[1][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[1][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[1][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[1][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[1][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[1][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[1][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[1][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[1][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[1][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[1][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[1][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[1][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[1][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[1][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[1][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[1][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[1][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[1][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[1][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[1][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[1][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[1][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[1][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[1][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[1][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[1][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[1][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[1][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[1][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[1][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[1][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[1][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[1][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[1][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[1][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[1][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[1][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[1][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[1][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[1][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[1][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[1][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[1][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[1][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[1][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[1][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[1][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[1][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[1][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[1][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[1][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[1][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[1][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[1][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[1][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[1][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[1][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[1][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[1][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[1][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[1][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[1][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[1][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[1][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[1][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[1][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[1][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[1][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[1][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[1][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[1][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[1][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[1][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[1][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[1][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[1][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[1][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[1][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[1][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[1][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[1][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[1][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[1][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[1][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[1][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[1][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[1][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[1][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[1][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[1][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[1][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[1][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[1][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[1][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[1][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[1][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[1][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[1][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[1][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[1][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[1][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[1][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[1][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[1][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[1][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[1][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[1][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[1][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[1][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[1][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[1][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[1][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[1][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[1][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[1][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[1][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[1][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[1][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[1][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[1][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[1][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[1][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[1][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[1][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[1][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[1][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[1][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[1][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[1][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[1][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[1][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[1][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[1][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[1][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[1][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[1][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[1][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[1][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[1][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[1][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[1][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[1][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[1][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[1][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[1][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[1][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[1][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[1][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[1][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[1][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[1][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[1][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[1][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[1][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[1][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[1][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[1][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[1][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[1][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 1, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[1][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[1][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[1][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[1][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[1][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[1].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[1][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[2][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[2][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[2][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[2][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[2][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[2][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[2][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[2][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[2][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[2][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[2][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[2][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[2][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[2][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[2][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[2][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[2][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[2][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[2][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[2][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[2][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[2][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[2][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[2][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[2][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[2][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[2][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[2][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[2][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[2][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[2][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[2][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[2][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[2][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[2][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[2][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[2][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[2][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[2][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[2][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[2][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[2][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[2][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[2][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[2][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[2][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[2][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[2][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[2][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[2][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[2][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[2][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[2][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[2][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[2][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[2][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[2][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[2][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[2][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[2][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[2][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[2][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[2][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[2][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[2][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[2][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[2][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[2][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[2][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[2][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[2][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[2][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[2][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[2][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[2][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[2][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[2][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[2][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[2][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[2][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[2][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[2][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[2][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[2][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[2][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[2][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[2][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[2][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[2][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[2][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[2][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[2][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[2][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[2][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[2][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[2][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[2][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[2][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[2][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[2][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[2][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[2][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[2][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[2][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[2][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[2][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[2][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[2][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[2][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[2][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[2][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[2][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[2][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[2][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[2][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[2][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[2][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[2][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[2][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[2][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[2][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[2][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[2][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[2][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[2][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[2][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[2][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[2][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[2][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[2][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[2][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[2][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[2][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[2][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[2][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[2][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[2][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[2][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[2][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[2][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[2][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[2][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[2][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[2][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[2][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[2][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[2][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[2][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[2][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[2][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[2][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[2][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[2][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[2][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[2][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[2][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[2][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[2][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[2][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[2][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[2][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[2][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[2][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[2][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[2][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[2][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[2][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[2][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[2][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[2][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[2][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[2][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[2][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[2][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[2][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[2][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[2][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[2][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[2][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[2][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[2][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[2][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[2][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[2][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[2][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[2][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 2, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[2][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[2][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[2][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[2][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[2][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[2].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[2][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[3][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[3][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[3][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[3][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[3][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[3][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[3][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[3][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[3][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[3][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[3][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[3][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[3][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[3][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[3][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[3][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[3][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[3][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[3][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[3][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[3][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[3][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[3][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[3][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[3][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[3][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[3][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[3][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[3][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[3][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[3][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[3][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[3][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[3][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[3][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[3][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[3][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[3][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[3][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[3][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[3][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[3][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[3][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[3][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[3][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[3][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[3][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[3][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[3][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[3][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[3][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[3][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[3][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[3][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[3][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[3][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[3][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[3][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[3][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[3][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[3][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[3][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[3][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[3][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[3][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[3][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[3][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[3][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[3][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[3][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[3][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[3][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[3][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[3][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[3][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[3][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[3][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[3][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[3][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[3][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[3][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[3][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[3][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[3][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[3][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[3][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[3][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[3][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[3][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[3][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[3][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[3][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[3][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[3][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[3][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[3][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[3][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[3][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[3][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[3][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[3][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[3][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[3][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[3][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[3][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[3][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[3][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[3][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[3][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[3][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[3][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[3][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[3][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[3][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[3][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[3][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[3][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[3][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[3][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[3][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[3][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[3][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[3][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[3][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[3][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[3][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[3][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[3][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[3][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[3][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[3][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[3][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[3][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[3][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[3][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[3][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[3][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[3][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[3][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[3][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[3][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[3][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[3][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[3][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[3][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[3][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[3][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[3][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[3][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[3][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[3][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[3][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[3][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[3][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[3][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[3][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[3][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[3][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[3][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[3][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[3][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[3][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[3][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[3][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[3][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[3][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[3][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[3][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[3][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[3][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[3][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[3][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[3][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[3][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[3][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[3][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[3][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[3][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[3][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[3][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[3][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[3][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[3][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[3][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[3][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[3][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 3, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[3][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[3][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[3][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[3][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[3][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[3].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[3][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[4][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[4][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[4][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[4][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[4][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[4][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[4][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[4][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[4][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[4][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[4][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[4][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[4][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[4][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[4][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[4][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[4][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[4][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[4][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[4][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[4][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[4][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[4][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[4][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[4][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[4][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[4][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[4][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[4][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[4][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[4][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[4][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[4][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[4][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[4][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[4][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[4][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[4][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[4][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[4][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[4][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[4][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[4][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[4][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[4][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[4][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[4][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[4][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[4][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[4][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[4][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[4][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[4][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[4][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[4][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[4][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[4][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[4][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[4][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[4][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[4][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[4][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[4][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[4][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[4][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[4][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[4][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[4][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[4][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[4][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[4][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[4][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[4][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[4][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[4][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[4][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[4][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[4][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[4][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[4][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[4][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[4][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[4][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[4][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[4][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[4][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[4][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[4][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[4][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[4][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[4][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[4][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[4][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[4][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[4][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[4][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[4][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[4][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[4][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[4][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[4][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[4][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[4][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[4][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[4][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[4][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[4][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[4][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[4][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[4][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[4][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[4][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[4][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[4][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[4][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[4][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[4][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[4][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[4][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[4][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[4][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[4][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[4][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[4][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[4][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[4][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[4][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[4][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[4][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[4][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[4][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[4][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[4][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[4][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[4][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[4][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[4][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[4][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[4][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[4][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[4][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[4][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[4][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[4][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[4][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[4][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[4][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[4][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[4][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[4][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[4][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[4][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[4][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[4][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[4][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[4][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[4][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[4][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[4][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[4][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[4][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[4][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[4][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[4][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[4][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[4][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[4][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[4][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[4][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[4][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[4][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[4][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[4][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[4][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[4][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[4][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[4][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[4][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[4][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[4][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[4][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[4][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[4][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[4][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[4][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[4][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 4, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[4][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[4][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[4][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[4][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[4][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[4].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[4][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[5][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[5][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[5][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[5][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[5][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[5][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[5][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[5][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[5][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[5][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[5][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[5][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[5][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[5][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[5][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[5][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[5][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[5][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[5][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[5][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[5][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[5][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[5][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[5][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[5][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[5][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[5][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[5][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[5][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[5][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[5][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[5][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[5][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[5][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[5][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[5][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[5][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[5][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[5][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[5][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[5][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[5][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[5][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[5][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[5][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[5][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[5][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[5][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[5][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[5][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[5][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[5][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[5][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[5][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[5][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[5][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[5][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[5][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[5][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[5][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[5][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[5][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[5][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[5][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[5][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[5][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[5][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[5][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[5][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[5][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[5][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[5][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[5][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[5][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[5][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[5][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[5][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[5][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[5][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[5][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[5][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[5][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[5][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[5][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[5][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[5][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[5][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[5][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[5][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[5][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[5][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[5][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[5][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[5][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[5][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[5][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[5][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[5][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[5][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[5][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[5][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[5][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[5][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[5][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[5][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[5][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[5][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[5][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[5][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[5][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[5][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[5][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[5][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[5][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[5][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[5][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[5][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[5][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[5][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[5][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[5][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[5][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[5][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[5][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[5][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[5][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[5][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[5][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[5][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[5][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[5][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[5][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[5][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[5][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[5][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[5][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[5][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[5][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[5][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[5][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[5][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[5][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[5][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[5][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[5][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[5][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[5][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[5][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[5][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[5][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[5][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[5][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[5][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[5][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[5][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[5][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[5][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[5][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[5][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[5][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[5][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[5][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[5][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[5][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[5][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[5][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[5][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[5][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[5][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[5][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[5][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[5][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[5][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[5][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[5][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[5][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[5][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[5][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[5][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[5][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[5][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[5][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[5][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[5][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[5][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[5][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 5, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[5][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[5][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[5][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[5][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[5][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[5].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[5][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[6][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[6][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[6][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[6][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[6][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[6][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[6][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[6][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[6][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[6][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[6][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[6][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[6][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[6][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[6][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[6][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[6][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[6][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[6][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[6][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[6][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[6][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[6][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[6][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[6][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[6][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[6][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[6][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[6][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[6][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[6][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[6][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[6][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[6][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[6][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[6][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[6][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[6][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[6][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[6][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[6][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[6][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[6][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[6][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[6][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[6][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[6][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[6][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[6][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[6][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[6][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[6][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[6][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[6][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[6][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[6][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[6][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[6][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[6][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[6][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[6][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[6][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[6][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[6][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[6][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[6][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[6][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[6][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[6][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[6][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[6][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[6][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[6][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[6][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[6][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[6][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[6][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[6][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[6][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[6][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[6][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[6][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[6][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[6][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[6][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[6][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[6][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[6][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[6][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[6][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[6][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[6][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[6][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[6][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[6][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[6][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[6][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[6][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[6][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[6][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[6][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[6][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[6][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[6][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[6][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[6][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[6][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[6][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[6][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[6][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[6][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[6][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[6][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[6][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[6][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[6][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[6][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[6][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[6][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[6][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[6][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[6][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[6][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[6][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[6][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[6][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[6][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[6][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[6][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[6][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[6][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[6][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[6][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[6][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[6][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[6][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[6][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[6][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[6][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[6][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[6][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[6][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[6][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[6][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[6][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[6][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[6][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[6][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[6][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[6][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[6][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[6][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[6][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[6][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[6][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[6][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[6][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[6][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[6][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[6][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[6][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[6][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[6][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[6][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[6][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[6][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[6][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[6][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[6][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[6][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[6][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[6][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[6][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[6][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[6][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[6][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[6][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[6][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[6][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[6][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[6][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[6][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[6][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[6][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[6][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[6][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 6, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[6][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[6][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[6][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[6][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[6][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[6].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[6][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[7][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[7][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[7][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[7][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[7][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[7][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[7][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[7][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[7][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[7][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[7][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[7][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[7][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[7][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[7][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[7][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[7][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[7][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[7][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[7][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[7][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[7][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[7][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[7][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[7][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[7][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[7][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[7][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[7][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[7][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[7][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[7][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[7][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[7][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[7][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[7][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[7][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[7][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[7][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[7][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[7][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[7][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[7][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[7][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[7][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[7][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[7][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[7][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[7][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[7][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[7][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[7][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[7][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[7][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[7][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[7][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[7][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[7][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[7][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[7][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[7][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[7][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[7][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[7][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[7][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[7][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[7][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[7][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[7][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[7][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[7][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[7][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[7][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[7][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[7][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[7][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[7][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[7][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[7][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[7][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[7][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[7][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[7][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[7][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[7][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[7][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[7][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[7][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[7][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[7][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[7][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[7][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[7][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[7][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[7][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[7][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[7][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[7][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[7][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[7][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[7][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[7][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[7][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[7][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[7][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[7][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[7][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[7][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[7][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[7][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[7][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[7][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[7][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[7][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[7][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[7][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[7][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[7][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[7][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[7][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[7][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[7][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[7][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[7][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[7][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[7][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[7][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[7][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[7][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[7][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[7][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[7][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[7][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[7][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[7][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[7][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[7][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[7][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[7][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[7][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[7][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[7][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[7][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[7][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[7][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[7][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[7][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[7][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[7][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[7][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[7][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[7][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[7][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[7][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[7][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[7][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[7][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[7][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[7][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[7][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[7][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[7][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[7][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[7][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[7][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[7][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[7][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[7][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[7][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[7][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[7][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[7][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[7][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[7][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[7][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[7][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[7][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[7][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[7][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[7][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[7][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[7][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[7][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[7][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[7][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[7][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 7, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[7][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[7][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[7][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[7][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[7][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[7].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[7][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[8][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[8][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[8][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[8][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[8][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[8][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[8][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[8][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[8][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[8][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[8][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[8][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[8][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[8][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[8][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[8][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[8][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[8][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[8][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[8][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[8][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[8][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[8][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[8][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[8][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[8][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[8][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[8][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[8][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[8][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[8][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[8][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[8][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[8][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[8][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[8][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[8][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[8][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[8][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[8][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[8][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[8][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[8][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[8][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[8][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[8][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[8][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[8][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[8][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[8][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[8][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[8][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[8][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[8][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[8][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[8][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[8][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[8][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[8][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[8][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[8][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[8][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[8][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[8][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[8][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[8][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[8][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[8][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[8][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[8][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[8][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[8][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[8][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[8][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[8][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[8][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[8][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[8][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[8][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[8][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[8][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[8][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[8][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[8][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[8][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[8][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[8][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[8][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[8][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[8][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[8][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[8][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[8][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[8][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[8][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[8][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[8][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[8][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[8][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[8][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[8][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[8][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[8][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[8][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[8][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[8][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[8][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[8][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[8][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[8][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[8][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[8][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[8][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[8][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[8][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[8][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[8][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[8][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[8][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[8][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[8][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[8][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[8][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[8][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[8][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[8][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[8][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[8][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[8][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[8][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[8][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[8][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[8][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[8][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[8][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[8][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[8][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[8][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[8][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[8][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[8][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[8][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[8][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[8][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[8][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[8][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[8][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[8][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[8][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[8][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[8][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[8][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[8][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[8][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[8][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[8][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[8][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[8][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[8][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[8][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[8][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[8][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[8][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[8][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[8][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[8][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[8][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[8][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[8][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[8][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[8][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[8][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[8][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[8][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[8][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[8][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[8][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[8][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[8][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[8][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[8][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[8][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[8][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[8][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[8][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[8][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 8, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[8][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[8][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[8][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[8][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[8][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[8].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[8][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[9][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[9][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[9][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[9][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[9][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[9][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[9][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[9][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[9][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[9][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[9][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[9][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[9][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[9][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[9][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[9][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[9][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[9][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[9][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[9][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[9][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[9][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[9][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[9][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[9][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[9][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[9][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[9][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[9][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[9][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[9][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[9][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[9][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[9][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[9][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[9][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[9][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[9][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[9][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[9][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[9][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[9][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[9][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[9][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[9][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[9][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[9][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[9][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[9][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[9][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[9][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[9][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[9][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[9][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[9][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[9][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[9][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[9][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[9][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[9][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[9][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[9][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[9][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[9][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[9][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[9][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[9][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[9][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[9][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[9][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[9][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[9][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[9][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[9][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[9][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[9][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[9][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[9][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[9][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[9][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[9][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[9][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[9][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[9][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[9][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[9][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[9][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[9][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[9][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[9][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[9][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[9][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[9][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[9][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[9][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[9][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[9][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[9][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[9][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[9][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[9][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[9][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[9][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[9][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[9][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[9][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[9][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[9][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[9][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[9][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[9][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[9][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[9][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[9][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[9][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[9][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[9][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[9][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[9][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[9][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[9][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[9][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[9][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[9][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[9][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[9][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[9][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[9][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[9][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[9][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[9][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[9][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[9][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[9][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[9][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[9][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[9][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[9][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[9][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[9][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[9][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[9][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[9][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[9][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[9][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[9][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[9][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[9][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[9][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[9][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[9][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[9][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[9][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[9][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[9][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[9][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[9][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[9][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[9][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[9][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[9][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[9][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[9][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[9][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[9][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[9][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[9][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[9][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[9][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[9][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[9][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[9][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[9][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[9][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[9][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[9][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[9][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[9][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[9][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[9][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[9][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[9][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[9][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[9][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[9][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[9][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 9, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[9][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[9][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[9][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[9][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[9][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[9].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[9][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[10][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[10][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[10][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[10][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[10][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[10][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[10][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[10][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[10][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[10][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[10][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[10][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[10][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[10][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[10][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[10][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[10][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[10][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[10][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[10][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[10][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[10][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[10][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[10][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[10][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[10][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[10][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[10][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[10][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[10][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[10][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[10][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[10][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[10][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[10][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[10][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[10][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[10][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[10][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[10][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[10][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[10][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[10][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[10][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[10][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[10][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[10][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[10][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[10][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[10][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[10][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[10][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[10][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[10][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[10][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[10][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[10][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[10][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[10][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[10][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[10][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[10][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[10][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[10][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[10][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[10][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[10][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[10][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[10][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[10][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[10][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[10][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[10][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[10][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[10][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[10][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[10][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[10][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[10][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[10][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[10][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[10][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[10][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[10][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[10][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[10][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[10][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[10][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[10][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[10][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[10][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[10][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[10][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[10][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[10][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[10][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[10][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[10][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[10][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[10][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[10][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[10][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[10][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[10][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[10][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[10][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[10][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[10][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[10][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[10][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[10][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[10][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[10][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[10][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[10][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[10][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[10][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[10][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[10][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[10][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[10][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[10][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[10][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[10][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[10][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[10][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[10][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[10][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[10][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[10][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[10][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[10][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[10][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[10][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[10][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[10][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[10][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[10][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[10][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[10][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[10][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[10][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[10][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[10][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[10][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[10][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[10][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[10][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[10][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[10][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[10][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[10][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[10][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[10][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[10][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[10][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[10][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[10][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[10][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[10][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[10][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[10][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[10][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[10][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[10][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[10][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[10][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[10][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[10][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[10][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[10][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[10][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[10][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[10][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[10][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[10][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[10][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[10][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[10][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[10][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[10][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[10][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[10][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[10][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[10][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[10][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 10, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[10][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[10][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[10][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[10][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[10][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[10].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[10][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[11][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[11][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[11][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[11][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[11][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[11][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[11][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[11][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[11][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[11][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[11][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[11][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[11][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[11][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[11][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[11][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[11][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[11][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[11][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[11][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[11][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[11][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[11][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[11][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[11][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[11][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[11][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[11][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[11][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[11][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[11][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[11][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[11][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[11][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[11][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[11][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[11][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[11][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[11][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[11][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[11][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[11][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[11][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[11][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[11][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[11][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[11][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[11][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[11][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[11][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[11][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[11][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[11][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[11][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[11][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[11][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[11][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[11][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[11][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[11][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[11][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[11][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[11][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[11][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[11][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[11][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[11][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[11][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[11][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[11][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[11][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[11][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[11][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[11][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[11][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[11][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[11][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[11][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[11][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[11][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[11][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[11][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[11][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[11][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[11][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[11][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[11][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[11][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[11][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[11][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[11][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[11][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[11][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[11][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[11][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[11][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[11][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[11][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[11][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[11][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[11][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[11][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[11][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[11][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[11][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[11][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[11][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[11][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[11][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[11][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[11][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[11][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[11][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[11][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[11][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[11][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[11][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[11][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[11][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[11][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[11][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[11][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[11][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[11][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[11][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[11][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[11][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[11][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[11][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[11][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[11][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[11][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[11][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[11][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[11][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[11][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[11][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[11][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[11][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[11][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[11][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[11][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[11][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[11][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[11][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[11][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[11][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[11][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[11][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[11][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[11][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[11][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[11][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[11][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[11][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[11][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[11][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[11][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[11][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[11][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[11][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[11][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[11][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[11][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[11][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[11][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[11][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[11][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[11][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[11][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[11][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[11][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[11][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[11][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[11][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[11][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[11][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[11][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[11][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[11][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[11][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[11][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[11][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[11][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[11][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[11][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 11, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[11][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[11][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[11][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[11][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[11][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[11].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[11][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[12][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[12][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[12][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[12][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[12][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[12][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[12][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[12][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[12][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[12][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[12][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[12][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[12][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[12][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[12][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[12][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[12][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[12][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[12][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[12][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[12][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[12][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[12][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[12][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[12][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[12][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[12][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[12][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[12][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[12][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[12][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[12][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[12][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[12][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[12][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[12][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[12][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[12][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[12][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[12][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[12][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[12][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[12][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[12][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[12][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[12][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[12][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[12][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[12][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[12][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[12][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[12][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[12][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[12][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[12][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[12][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[12][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[12][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[12][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[12][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[12][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[12][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[12][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[12][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[12][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[12][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[12][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[12][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[12][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[12][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[12][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[12][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[12][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[12][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[12][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[12][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[12][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[12][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[12][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[12][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[12][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[12][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[12][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[12][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[12][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[12][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[12][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[12][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[12][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[12][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[12][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[12][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[12][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[12][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[12][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[12][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[12][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[12][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[12][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[12][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[12][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[12][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[12][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[12][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[12][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[12][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[12][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[12][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[12][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[12][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[12][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[12][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[12][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[12][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[12][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[12][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[12][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[12][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[12][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[12][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[12][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[12][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[12][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[12][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[12][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[12][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[12][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[12][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[12][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[12][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[12][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[12][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[12][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[12][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[12][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[12][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[12][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[12][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[12][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[12][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[12][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[12][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[12][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[12][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[12][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[12][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[12][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[12][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[12][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[12][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[12][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[12][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[12][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[12][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[12][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[12][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[12][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[12][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[12][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[12][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[12][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[12][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[12][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[12][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[12][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[12][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[12][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[12][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[12][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[12][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[12][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[12][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[12][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[12][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[12][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[12][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[12][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[12][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[12][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[12][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[12][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[12][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[12][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[12][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[12][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[12][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 12, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[12][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[12][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[12][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[12][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[12][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[12].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[12][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[13][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[13][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[13][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[13][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[13][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[13][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[13][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[13][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[13][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[13][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[13][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[13][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[13][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[13][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[13][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[13][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[13][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[13][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[13][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[13][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[13][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[13][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[13][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[13][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[13][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[13][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[13][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[13][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[13][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[13][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[13][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[13][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[13][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[13][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[13][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[13][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[13][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[13][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[13][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[13][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[13][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[13][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[13][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[13][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[13][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[13][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[13][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[13][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[13][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[13][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[13][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[13][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[13][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[13][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[13][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[13][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[13][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[13][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[13][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[13][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[13][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[13][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[13][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[13][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[13][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[13][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[13][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[13][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[13][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[13][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[13][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[13][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[13][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[13][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[13][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[13][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[13][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[13][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[13][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[13][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[13][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[13][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[13][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[13][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[13][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[13][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[13][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[13][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[13][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[13][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[13][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[13][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[13][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[13][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[13][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[13][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[13][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[13][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[13][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[13][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[13][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[13][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[13][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[13][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[13][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[13][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[13][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[13][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[13][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[13][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[13][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[13][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[13][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[13][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[13][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[13][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[13][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[13][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[13][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[13][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[13][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[13][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[13][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[13][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[13][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[13][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[13][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[13][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[13][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[13][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[13][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[13][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[13][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[13][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[13][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[13][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[13][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[13][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[13][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[13][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[13][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[13][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[13][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[13][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[13][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[13][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[13][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[13][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[13][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[13][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[13][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[13][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[13][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[13][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[13][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[13][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[13][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[13][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[13][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[13][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[13][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[13][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[13][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[13][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[13][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[13][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[13][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[13][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[13][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[13][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[13][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[13][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[13][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[13][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[13][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[13][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[13][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[13][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[13][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[13][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[13][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[13][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[13][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[13][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[13][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[13][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 13, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[13][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[13][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[13][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[13][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[13][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[13].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[13][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[14][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[14][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[14][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[14][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[14][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[14][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[14][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[14][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[14][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[14][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[14][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[14][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[14][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[14][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[14][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[14][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[14][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[14][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[14][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[14][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[14][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[14][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[14][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[14][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[14][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[14][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[14][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[14][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[14][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[14][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[14][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[14][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[14][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[14][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[14][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[14][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[14][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[14][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[14][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[14][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[14][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[14][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[14][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[14][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[14][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[14][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[14][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[14][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[14][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[14][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[14][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[14][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[14][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[14][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[14][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[14][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[14][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[14][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[14][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[14][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[14][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[14][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[14][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[14][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[14][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[14][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[14][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[14][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[14][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[14][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[14][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[14][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[14][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[14][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[14][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[14][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[14][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[14][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[14][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[14][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[14][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[14][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[14][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[14][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[14][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[14][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[14][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[14][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[14][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[14][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[14][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[14][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[14][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[14][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[14][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[14][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[14][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[14][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[14][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[14][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[14][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[14][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[14][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[14][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[14][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[14][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[14][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[14][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[14][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[14][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[14][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[14][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[14][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[14][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[14][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[14][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[14][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[14][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[14][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[14][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[14][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[14][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[14][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[14][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[14][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[14][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[14][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[14][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[14][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[14][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[14][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[14][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[14][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[14][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[14][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[14][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[14][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[14][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[14][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[14][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[14][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[14][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[14][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[14][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[14][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[14][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[14][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[14][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[14][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[14][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[14][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[14][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[14][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[14][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[14][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[14][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[14][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[14][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[14][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[14][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[14][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[14][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[14][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[14][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[14][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[14][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[14][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[14][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[14][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[14][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[14][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[14][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[14][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[14][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[14][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[14][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[14][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[14][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[14][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[14][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[14][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[14][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[14][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[14][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[14][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[14][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 14, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[14][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[14][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[14][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[14][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[14][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[14].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[14][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[15][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[15][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[15][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[15][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[15][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[15][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[15][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[15][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[15][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[15][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[15][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[15][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[15][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[15][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[15][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[15][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[15][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[15][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[15][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[15][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[15][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[15][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[15][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[15][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[15][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[15][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[15][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[15][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[15][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[15][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[15][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[15][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[15][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[15][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[15][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[15][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[15][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[15][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[15][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[15][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[15][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[15][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[15][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[15][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[15][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[15][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[15][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[15][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[15][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[15][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[15][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[15][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[15][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[15][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[15][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[15][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[15][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[15][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[15][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[15][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[15][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[15][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[15][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[15][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[15][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[15][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[15][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[15][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[15][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[15][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[15][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[15][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[15][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[15][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[15][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[15][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[15][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[15][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[15][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[15][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[15][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[15][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[15][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[15][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[15][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[15][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[15][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[15][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[15][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[15][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[15][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[15][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[15][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[15][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[15][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[15][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[15][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[15][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[15][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[15][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[15][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[15][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[15][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[15][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[15][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[15][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[15][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[15][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[15][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[15][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[15][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[15][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[15][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[15][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[15][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[15][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[15][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[15][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[15][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[15][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[15][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[15][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[15][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[15][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[15][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[15][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[15][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[15][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[15][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[15][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[15][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[15][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[15][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[15][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[15][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[15][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[15][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[15][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[15][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[15][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[15][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[15][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[15][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[15][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[15][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[15][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[15][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[15][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[15][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[15][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[15][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[15][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[15][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[15][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[15][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[15][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[15][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[15][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[15][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[15][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[15][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[15][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[15][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[15][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[15][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[15][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[15][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[15][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[15][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[15][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[15][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[15][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[15][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[15][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[15][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[15][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[15][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[15][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[15][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[15][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[15][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[15][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[15][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[15][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[15][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[15][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 15, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[15][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[15][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[15][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[15][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[15][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[15].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[15][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[16][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[16][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[16][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[16][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[16][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[16][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[16][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[16][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[16][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[16][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[16][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[16][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[16][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[16][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[16][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[16][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[16][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[16][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[16][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[16][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[16][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[16][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[16][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[16][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[16][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[16][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[16][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[16][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[16][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[16][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[16][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[16][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[16][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[16][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[16][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[16][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[16][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[16][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[16][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[16][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[16][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[16][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[16][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[16][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[16][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[16][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[16][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[16][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[16][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[16][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[16][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[16][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[16][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[16][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[16][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[16][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[16][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[16][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[16][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[16][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[16][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[16][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[16][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[16][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[16][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[16][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[16][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[16][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[16][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[16][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[16][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[16][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[16][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[16][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[16][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[16][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[16][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[16][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[16][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[16][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[16][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[16][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[16][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[16][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[16][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[16][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[16][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[16][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[16][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[16][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[16][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[16][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[16][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[16][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[16][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[16][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[16][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[16][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[16][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[16][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[16][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[16][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[16][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[16][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[16][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[16][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[16][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[16][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[16][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[16][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[16][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[16][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[16][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[16][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[16][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[16][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[16][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[16][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[16][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[16][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[16][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[16][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[16][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[16][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[16][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[16][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[16][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[16][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[16][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[16][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[16][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[16][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[16][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[16][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[16][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[16][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[16][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[16][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[16][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[16][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[16][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[16][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[16][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[16][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[16][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[16][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[16][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[16][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[16][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[16][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[16][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[16][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[16][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[16][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[16][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[16][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[16][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[16][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[16][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[16][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[16][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[16][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[16][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[16][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[16][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[16][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[16][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[16][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[16][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[16][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[16][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[16][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[16][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[16][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[16][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[16][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[16][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[16][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[16][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[16][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[16][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[16][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[16][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[16][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[16][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[16][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 16, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[16][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[16][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[16][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[16][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[16][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[16].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[16][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[17][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[17][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[17][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[17][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[17][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[17][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[17][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[17][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[17][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[17][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[17][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[17][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[17][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[17][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[17][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[17][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[17][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[17][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[17][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[17][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[17][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[17][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[17][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[17][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[17][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[17][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[17][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[17][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[17][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[17][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[17][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[17][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[17][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[17][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[17][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[17][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[17][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[17][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[17][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[17][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[17][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[17][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[17][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[17][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[17][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[17][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[17][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[17][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[17][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[17][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[17][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[17][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[17][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[17][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[17][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[17][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[17][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[17][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[17][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[17][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[17][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[17][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[17][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[17][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[17][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[17][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[17][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[17][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[17][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[17][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[17][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[17][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[17][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[17][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[17][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[17][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[17][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[17][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[17][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[17][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[17][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[17][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[17][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[17][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[17][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[17][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[17][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[17][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[17][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[17][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[17][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[17][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[17][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[17][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[17][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[17][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[17][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[17][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[17][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[17][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[17][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[17][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[17][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[17][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[17][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[17][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[17][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[17][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[17][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[17][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[17][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[17][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[17][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[17][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[17][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[17][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[17][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[17][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[17][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[17][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[17][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[17][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[17][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[17][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[17][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[17][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[17][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[17][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[17][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[17][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[17][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[17][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[17][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[17][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[17][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[17][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[17][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[17][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[17][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[17][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[17][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[17][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[17][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[17][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[17][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[17][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[17][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[17][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[17][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[17][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[17][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[17][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[17][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[17][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[17][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[17][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[17][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[17][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[17][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[17][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[17][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[17][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[17][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[17][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[17][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[17][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[17][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[17][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[17][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[17][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[17][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[17][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[17][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[17][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[17][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[17][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[17][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[17][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[17][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[17][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[17][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[17][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[17][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[17][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[17][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[17][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 17, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[17][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[17][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[17][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[17][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[17][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[17].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[17][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[18][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[18][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[18][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[18][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[18][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[18][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[18][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[18][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[18][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[18][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[18][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[18][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[18][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[18][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[18][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[18][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[18][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[18][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[18][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[18][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[18][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[18][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[18][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[18][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[18][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[18][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[18][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[18][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[18][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[18][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[18][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[18][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[18][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[18][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[18][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[18][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[18][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[18][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[18][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[18][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[18][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[18][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[18][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[18][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[18][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[18][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[18][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[18][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[18][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[18][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[18][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[18][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[18][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[18][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[18][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[18][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[18][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[18][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[18][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[18][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[18][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[18][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[18][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[18][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[18][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[18][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[18][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[18][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[18][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[18][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[18][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[18][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[18][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[18][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[18][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[18][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[18][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[18][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[18][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[18][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[18][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[18][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[18][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[18][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[18][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[18][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[18][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[18][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[18][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[18][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[18][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[18][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[18][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[18][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[18][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[18][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[18][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[18][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[18][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[18][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[18][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[18][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[18][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[18][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[18][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[18][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[18][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[18][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[18][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[18][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[18][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[18][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[18][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[18][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[18][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[18][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[18][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[18][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[18][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[18][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[18][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[18][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[18][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[18][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[18][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[18][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[18][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[18][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[18][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[18][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[18][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[18][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[18][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[18][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[18][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[18][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[18][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[18][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[18][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[18][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[18][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[18][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[18][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[18][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[18][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[18][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[18][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[18][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[18][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[18][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[18][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[18][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[18][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[18][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[18][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[18][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[18][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[18][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[18][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[18][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[18][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[18][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[18][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[18][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[18][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[18][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[18][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[18][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[18][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[18][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[18][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[18][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[18][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[18][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[18][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[18][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[18][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[18][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[18][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[18][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[18][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[18][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[18][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[18][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[18][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[18][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 18, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[18][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[18][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[18][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[18][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[18][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[18].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[18][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[19][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[19][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[19][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[19][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[19][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[19][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[19][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[19][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[19][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[19][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[19][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[19][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[19][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[19][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[19][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[19][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[19][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[19][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[19][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[19][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[19][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[19][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[19][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[19][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[19][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[19][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[19][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[19][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[19][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[19][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[19][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[19][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[19][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[19][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[19][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[19][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[19][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[19][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[19][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[19][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[19][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[19][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[19][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[19][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[19][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[19][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[19][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[19][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[19][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[19][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[19][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[19][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[19][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[19][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[19][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[19][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[19][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[19][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[19][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[19][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[19][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[19][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[19][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[19][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[19][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[19][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[19][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[19][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[19][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[19][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[19][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[19][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[19][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[19][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[19][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[19][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[19][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[19][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[19][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[19][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[19][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[19][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[19][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[19][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[19][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[19][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[19][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[19][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[19][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[19][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[19][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[19][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[19][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[19][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[19][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[19][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[19][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[19][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[19][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[19][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[19][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[19][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[19][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[19][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[19][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[19][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[19][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[19][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[19][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[19][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[19][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[19][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[19][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[19][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[19][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[19][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[19][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[19][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[19][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[19][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[19][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[19][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[19][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[19][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[19][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[19][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[19][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[19][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[19][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[19][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[19][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[19][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[19][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[19][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[19][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[19][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[19][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[19][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[19][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[19][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[19][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[19][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[19][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[19][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[19][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[19][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[19][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[19][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[19][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[19][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[19][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[19][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[19][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[19][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[19][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[19][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[19][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[19][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[19][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[19][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[19][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[19][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[19][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[19][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[19][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[19][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[19][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[19][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[19][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[19][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[19][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[19][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[19][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[19][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[19][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[19][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[19][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[19][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[19][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[19][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[19][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[19][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[19][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[19][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[19][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[19][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 19, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[19][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[19][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[19][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[19][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[19][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[19].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[19][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[20][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[20][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[20][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[20][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[20][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[20][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[20][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[20][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[20][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[20][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[20][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[20][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[20][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[20][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[20][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[20][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[20][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[20][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[20][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[20][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[20][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[20][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[20][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[20][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[20][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[20][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[20][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[20][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[20][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[20][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[20][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[20][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[20][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[20][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[20][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[20][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[20][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[20][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[20][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[20][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[20][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[20][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[20][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[20][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[20][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[20][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[20][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[20][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[20][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[20][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[20][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[20][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[20][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[20][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[20][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[20][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[20][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[20][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[20][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[20][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[20][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[20][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[20][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[20][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[20][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[20][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[20][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[20][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[20][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[20][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[20][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[20][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[20][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[20][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[20][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[20][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[20][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[20][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[20][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[20][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[20][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[20][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[20][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[20][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[20][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[20][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[20][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[20][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[20][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[20][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[20][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[20][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[20][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[20][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[20][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[20][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[20][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[20][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[20][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[20][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[20][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[20][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[20][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[20][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[20][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[20][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[20][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[20][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[20][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[20][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[20][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[20][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[20][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[20][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[20][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[20][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[20][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[20][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[20][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[20][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[20][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[20][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[20][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[20][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[20][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[20][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[20][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[20][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[20][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[20][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[20][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[20][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[20][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[20][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[20][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[20][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[20][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[20][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[20][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[20][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[20][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[20][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[20][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[20][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[20][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[20][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[20][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[20][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[20][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[20][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[20][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[20][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[20][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[20][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[20][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[20][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[20][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[20][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[20][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[20][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[20][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[20][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[20][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[20][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[20][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[20][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[20][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[20][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[20][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[20][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[20][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[20][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[20][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[20][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[20][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[20][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[20][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[20][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[20][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[20][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[20][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[20][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[20][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[20][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[20][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[20][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 20, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[20][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[20][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[20][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[20][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[20][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[20].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[20][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[21][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[21][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[21][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[21][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[21][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[21][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[21][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[21][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[21][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[21][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[21][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[21][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[21][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[21][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[21][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[21][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[21][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[21][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[21][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[21][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[21][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[21][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[21][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[21][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[21][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[21][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[21][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[21][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[21][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[21][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[21][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[21][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[21][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[21][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[21][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[21][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[21][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[21][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[21][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[21][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[21][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[21][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[21][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[21][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[21][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[21][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[21][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[21][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[21][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[21][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[21][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[21][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[21][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[21][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[21][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[21][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[21][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[21][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[21][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[21][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[21][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[21][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[21][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[21][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[21][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[21][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[21][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[21][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[21][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[21][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[21][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[21][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[21][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[21][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[21][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[21][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[21][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[21][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[21][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[21][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[21][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[21][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[21][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[21][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[21][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[21][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[21][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[21][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[21][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[21][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[21][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[21][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[21][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[21][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[21][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[21][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[21][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[21][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[21][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[21][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[21][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[21][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[21][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[21][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[21][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[21][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[21][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[21][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[21][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[21][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[21][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[21][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[21][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[21][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[21][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[21][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[21][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[21][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[21][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[21][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[21][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[21][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[21][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[21][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[21][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[21][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[21][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[21][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[21][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[21][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[21][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[21][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[21][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[21][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[21][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[21][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[21][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[21][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[21][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[21][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[21][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[21][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[21][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[21][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[21][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[21][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[21][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[21][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[21][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[21][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[21][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[21][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[21][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[21][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[21][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[21][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[21][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[21][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[21][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[21][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[21][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[21][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[21][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[21][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[21][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[21][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[21][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[21][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[21][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[21][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[21][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[21][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[21][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[21][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[21][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[21][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[21][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[21][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[21][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[21][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[21][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[21][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[21][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[21][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[21][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[21][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 21, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[21][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[21][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[21][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[21][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[21][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[21].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[21][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[22][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[22][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[22][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[22][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[22][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[22][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[22][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[22][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[22][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[22][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[22][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[22][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[22][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[22][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[22][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[22][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[22][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[22][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[22][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[22][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[22][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[22][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[22][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[22][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[22][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[22][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[22][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[22][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[22][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[22][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[22][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[22][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[22][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[22][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[22][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[22][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[22][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[22][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[22][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[22][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[22][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[22][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[22][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[22][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[22][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[22][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[22][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[22][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[22][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[22][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[22][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[22][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[22][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[22][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[22][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[22][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[22][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[22][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[22][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[22][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[22][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[22][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[22][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[22][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[22][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[22][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[22][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[22][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[22][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[22][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[22][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[22][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[22][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[22][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[22][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[22][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[22][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[22][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[22][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[22][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[22][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[22][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[22][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[22][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[22][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[22][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[22][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[22][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[22][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[22][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[22][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[22][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[22][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[22][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[22][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[22][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[22][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[22][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[22][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[22][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[22][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[22][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[22][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[22][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[22][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[22][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[22][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[22][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[22][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[22][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[22][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[22][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[22][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[22][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[22][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[22][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[22][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[22][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[22][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[22][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[22][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[22][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[22][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[22][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[22][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[22][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[22][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[22][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[22][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[22][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[22][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[22][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[22][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[22][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[22][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[22][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[22][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[22][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[22][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[22][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[22][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[22][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[22][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[22][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[22][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[22][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[22][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[22][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[22][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[22][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[22][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[22][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[22][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[22][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[22][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[22][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[22][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[22][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[22][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[22][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[22][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[22][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[22][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[22][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[22][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[22][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[22][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[22][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[22][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[22][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[22][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[22][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[22][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[22][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[22][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[22][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[22][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[22][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[22][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[22][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[22][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[22][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[22][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[22][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[22][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[22][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 22, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[22][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[22][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[22][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[22][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[22][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[22].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[22][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[23][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[23][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[23][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[23][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[23][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[23][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[23][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[23][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[23][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[23][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[23][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[23][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[23][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[23][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[23][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[23][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[23][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[23][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[23][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[23][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[23][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[23][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[23][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[23][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[23][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[23][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[23][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[23][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[23][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[23][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[23][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[23][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[23][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[23][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[23][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[23][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[23][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[23][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[23][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[23][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[23][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[23][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[23][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[23][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[23][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[23][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[23][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[23][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[23][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[23][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[23][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[23][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[23][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[23][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[23][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[23][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[23][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[23][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[23][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[23][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[23][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[23][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[23][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[23][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[23][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[23][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[23][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[23][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[23][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[23][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[23][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[23][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[23][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[23][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[23][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[23][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[23][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[23][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[23][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[23][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[23][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[23][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[23][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[23][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[23][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[23][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[23][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[23][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[23][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[23][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[23][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[23][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[23][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[23][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[23][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[23][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[23][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[23][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[23][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[23][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[23][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[23][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[23][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[23][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[23][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[23][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[23][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[23][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[23][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[23][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[23][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[23][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[23][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[23][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[23][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[23][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[23][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[23][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[23][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[23][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[23][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[23][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[23][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[23][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[23][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[23][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[23][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[23][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[23][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[23][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[23][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[23][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[23][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[23][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[23][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[23][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[23][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[23][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[23][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[23][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[23][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[23][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[23][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[23][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[23][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[23][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[23][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[23][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[23][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[23][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[23][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[23][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[23][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[23][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[23][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[23][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[23][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[23][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[23][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[23][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[23][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[23][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[23][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[23][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[23][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[23][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[23][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[23][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[23][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[23][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[23][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[23][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[23][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[23][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[23][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[23][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[23][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[23][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[23][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[23][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[23][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[23][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[23][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[23][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[23][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[23][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 23, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[23][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[23][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[23][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[23][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[23][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[23].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[23][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[24][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[24][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[24][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[24][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[24][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[24][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[24][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[24][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[24][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[24][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[24][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[24][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[24][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[24][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[24][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[24][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[24][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[24][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[24][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[24][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[24][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[24][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[24][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[24][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[24][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[24][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[24][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[24][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[24][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[24][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[24][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[24][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[24][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[24][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[24][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[24][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[24][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[24][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[24][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[24][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[24][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[24][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[24][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[24][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[24][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[24][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[24][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[24][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[24][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[24][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[24][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[24][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[24][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[24][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[24][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[24][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[24][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[24][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[24][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[24][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[24][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[24][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[24][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[24][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[24][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[24][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[24][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[24][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[24][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[24][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[24][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[24][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[24][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[24][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[24][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[24][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[24][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[24][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[24][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[24][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[24][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[24][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[24][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[24][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[24][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[24][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[24][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[24][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[24][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[24][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[24][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[24][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[24][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[24][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[24][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[24][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[24][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[24][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[24][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[24][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[24][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[24][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[24][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[24][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[24][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[24][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[24][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[24][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[24][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[24][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[24][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[24][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[24][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[24][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[24][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[24][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[24][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[24][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[24][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[24][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[24][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[24][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[24][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[24][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[24][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[24][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[24][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[24][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[24][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[24][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[24][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[24][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[24][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[24][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[24][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[24][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[24][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[24][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[24][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[24][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[24][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[24][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[24][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[24][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[24][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[24][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[24][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[24][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[24][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[24][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[24][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[24][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[24][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[24][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[24][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[24][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[24][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[24][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[24][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[24][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[24][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[24][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[24][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[24][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[24][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[24][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[24][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[24][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[24][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[24][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[24][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[24][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[24][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[24][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[24][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[24][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[24][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[24][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[24][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[24][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[24][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[24][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[24][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[24][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[24][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[24][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 24, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[24][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[24][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[24][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[24][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[24][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[24].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[24][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[25][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[25][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[25][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[25][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[25][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[25][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[25][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[25][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[25][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[25][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[25][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[25][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[25][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[25][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[25][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[25][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[25][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[25][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[25][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[25][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[25][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[25][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[25][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[25][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[25][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[25][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[25][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[25][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[25][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[25][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[25][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[25][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[25][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[25][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[25][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[25][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[25][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[25][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[25][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[25][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[25][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[25][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[25][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[25][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[25][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[25][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[25][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[25][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[25][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[25][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[25][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[25][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[25][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[25][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[25][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[25][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[25][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[25][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[25][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[25][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[25][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[25][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[25][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[25][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[25][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[25][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[25][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[25][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[25][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[25][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[25][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[25][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[25][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[25][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[25][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[25][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[25][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[25][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[25][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[25][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[25][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[25][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[25][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[25][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[25][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[25][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[25][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[25][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[25][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[25][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[25][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[25][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[25][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[25][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[25][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[25][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[25][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[25][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[25][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[25][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[25][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[25][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[25][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[25][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[25][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[25][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[25][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[25][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[25][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[25][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[25][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[25][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[25][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[25][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[25][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[25][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[25][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[25][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[25][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[25][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[25][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[25][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[25][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[25][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[25][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[25][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[25][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[25][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[25][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[25][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[25][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[25][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[25][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[25][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[25][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[25][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[25][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[25][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[25][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[25][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[25][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[25][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[25][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[25][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[25][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[25][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[25][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[25][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[25][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[25][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[25][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[25][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[25][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[25][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[25][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[25][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[25][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[25][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[25][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[25][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[25][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[25][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[25][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[25][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[25][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[25][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[25][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[25][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[25][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[25][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[25][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[25][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[25][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[25][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[25][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[25][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[25][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[25][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[25][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[25][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[25][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[25][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[25][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[25][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[25][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[25][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 25, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[25][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[25][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[25][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[25][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[25][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[25].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[25][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[26][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[26][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[26][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[26][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[26][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[26][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[26][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[26][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[26][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[26][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[26][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[26][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[26][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[26][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[26][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[26][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[26][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[26][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[26][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[26][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[26][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[26][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[26][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[26][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[26][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[26][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[26][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[26][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[26][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[26][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[26][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[26][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[26][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[26][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[26][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[26][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[26][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[26][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[26][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[26][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[26][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[26][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[26][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[26][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[26][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[26][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[26][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[26][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[26][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[26][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[26][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[26][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[26][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[26][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[26][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[26][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[26][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[26][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[26][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[26][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[26][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[26][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[26][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[26][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[26][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[26][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[26][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[26][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[26][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[26][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[26][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[26][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[26][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[26][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[26][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[26][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[26][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[26][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[26][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[26][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[26][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[26][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[26][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[26][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[26][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[26][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[26][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[26][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[26][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[26][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[26][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[26][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[26][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[26][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[26][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[26][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[26][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[26][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[26][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[26][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[26][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[26][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[26][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[26][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[26][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[26][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[26][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[26][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[26][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[26][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[26][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[26][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[26][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[26][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[26][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[26][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[26][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[26][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[26][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[26][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[26][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[26][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[26][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[26][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[26][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[26][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[26][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[26][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[26][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[26][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[26][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[26][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[26][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[26][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[26][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[26][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[26][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[26][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[26][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[26][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[26][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[26][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[26][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[26][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[26][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[26][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[26][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[26][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[26][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[26][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[26][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[26][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[26][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[26][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[26][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[26][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[26][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[26][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[26][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[26][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[26][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[26][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[26][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[26][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[26][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[26][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[26][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[26][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[26][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[26][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[26][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[26][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[26][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[26][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[26][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[26][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[26][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[26][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[26][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[26][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[26][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[26][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[26][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[26][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[26][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[26][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 26, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[26][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[26][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[26][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[26][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[26][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[26].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[26][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[27][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[27][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[27][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[27][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[27][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[27][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[27][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[27][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[27][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[27][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[27][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[27][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[27][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[27][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[27][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[27][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[27][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[27][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[27][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[27][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[27][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[27][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[27][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[27][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[27][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[27][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[27][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[27][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[27][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[27][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[27][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[27][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[27][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[27][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[27][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[27][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[27][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[27][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[27][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[27][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[27][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[27][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[27][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[27][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[27][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[27][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[27][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[27][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[27][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[27][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[27][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[27][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[27][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[27][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[27][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[27][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[27][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[27][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[27][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[27][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[27][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[27][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[27][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[27][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[27][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[27][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[27][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[27][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[27][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[27][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[27][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[27][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[27][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[27][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[27][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[27][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[27][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[27][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[27][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[27][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[27][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[27][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[27][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[27][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[27][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[27][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[27][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[27][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[27][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[27][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[27][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[27][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[27][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[27][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[27][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[27][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[27][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[27][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[27][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[27][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[27][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[27][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[27][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[27][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[27][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[27][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[27][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[27][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[27][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[27][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[27][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[27][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[27][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[27][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[27][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[27][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[27][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[27][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[27][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[27][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[27][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[27][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[27][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[27][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[27][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[27][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[27][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[27][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[27][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[27][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[27][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[27][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[27][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[27][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[27][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[27][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[27][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[27][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[27][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[27][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[27][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[27][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[27][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[27][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[27][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[27][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[27][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[27][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[27][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[27][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[27][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[27][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[27][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[27][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[27][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[27][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[27][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[27][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[27][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[27][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[27][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[27][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[27][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[27][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[27][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[27][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[27][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[27][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[27][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[27][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[27][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[27][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[27][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[27][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[27][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[27][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[27][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[27][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[27][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[27][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[27][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[27][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[27][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[27][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[27][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[27][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 27, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[27][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[27][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[27][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[27][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[27][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[27].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[27][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[28][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[28][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[28][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[28][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[28][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[28][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[28][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[28][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[28][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[28][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[28][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[28][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[28][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[28][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[28][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[28][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[28][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[28][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[28][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[28][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[28][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[28][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[28][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[28][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[28][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[28][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[28][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[28][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[28][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[28][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[28][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[28][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[28][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[28][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[28][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[28][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[28][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[28][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[28][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[28][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[28][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[28][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[28][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[28][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[28][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[28][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[28][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[28][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[28][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[28][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[28][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[28][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[28][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[28][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[28][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[28][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[28][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[28][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[28][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[28][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[28][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[28][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[28][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[28][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[28][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[28][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[28][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[28][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[28][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[28][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[28][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[28][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[28][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[28][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[28][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[28][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[28][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[28][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[28][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[28][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[28][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[28][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[28][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[28][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[28][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[28][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[28][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[28][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[28][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[28][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[28][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[28][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[28][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[28][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[28][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[28][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[28][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[28][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[28][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[28][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[28][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[28][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[28][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[28][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[28][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[28][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[28][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[28][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[28][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[28][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[28][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[28][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[28][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[28][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[28][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[28][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[28][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[28][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[28][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[28][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[28][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[28][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[28][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[28][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[28][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[28][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[28][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[28][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[28][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[28][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[28][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[28][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[28][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[28][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[28][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[28][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[28][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[28][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[28][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[28][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[28][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[28][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[28][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[28][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[28][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[28][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[28][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[28][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[28][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[28][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[28][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[28][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[28][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[28][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[28][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[28][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[28][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[28][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[28][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[28][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[28][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[28][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[28][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[28][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[28][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[28][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[28][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[28][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[28][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[28][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[28][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[28][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[28][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[28][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[28][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[28][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[28][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[28][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[28][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[28][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[28][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[28][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[28][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[28][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[28][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[28][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 28, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[28][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[28][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[28][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[28][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[28][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[28].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[28][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[29][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[29][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[29][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[29][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[29][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[29][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[29][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[29][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[29][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[29][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[29][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[29][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[29][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[29][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[29][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[29][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[29][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[29][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[29][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[29][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[29][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[29][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[29][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[29][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[29][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[29][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[29][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[29][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[29][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[29][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[29][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[29][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[29][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[29][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[29][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[29][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[29][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[29][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[29][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[29][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[29][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[29][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[29][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[29][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[29][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[29][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[29][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[29][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[29][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[29][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[29][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[29][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[29][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[29][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[29][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[29][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[29][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[29][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[29][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[29][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[29][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[29][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[29][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[29][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[29][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[29][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[29][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[29][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[29][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[29][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[29][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[29][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[29][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[29][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[29][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[29][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[29][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[29][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[29][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[29][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[29][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[29][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[29][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[29][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[29][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[29][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[29][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[29][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[29][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[29][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[29][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[29][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[29][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[29][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[29][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[29][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[29][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[29][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[29][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[29][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[29][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[29][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[29][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[29][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[29][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[29][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[29][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[29][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[29][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[29][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[29][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[29][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[29][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[29][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[29][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[29][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[29][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[29][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[29][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[29][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[29][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[29][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[29][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[29][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[29][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[29][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[29][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[29][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[29][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[29][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[29][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[29][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[29][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[29][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[29][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[29][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[29][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[29][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[29][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[29][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[29][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[29][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[29][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[29][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[29][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[29][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[29][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[29][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[29][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[29][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[29][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[29][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[29][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[29][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[29][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[29][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[29][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[29][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[29][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[29][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[29][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[29][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[29][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[29][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[29][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[29][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[29][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[29][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[29][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[29][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[29][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[29][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[29][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[29][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[29][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[29][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[29][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[29][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[29][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[29][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[29][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[29][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[29][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[29][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[29][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[29][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 29, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[29][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[29][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[29][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[29][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[29][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[29].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[29][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[30][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[30][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[30][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[30][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[30][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[30][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[30][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[30][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[30][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[30][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[30][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[30][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[30][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[30][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[30][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[30][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[30][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[30][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[30][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[30][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[30][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[30][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[30][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[30][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[30][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[30][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[30][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[30][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[30][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[30][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[30][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[30][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[30][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[30][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[30][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[30][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[30][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[30][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[30][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[30][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[30][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[30][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[30][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[30][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[30][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[30][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[30][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[30][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[30][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[30][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[30][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[30][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[30][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[30][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[30][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[30][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[30][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[30][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[30][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[30][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[30][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[30][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[30][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[30][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[30][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[30][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[30][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[30][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[30][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[30][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[30][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[30][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[30][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[30][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[30][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[30][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[30][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[30][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[30][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[30][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[30][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[30][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[30][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[30][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[30][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[30][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[30][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[30][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[30][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[30][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[30][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[30][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[30][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[30][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[30][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[30][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[30][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[30][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[30][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[30][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[30][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[30][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[30][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[30][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[30][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[30][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[30][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[30][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[30][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[30][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[30][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[30][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[30][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[30][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[30][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[30][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[30][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[30][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[30][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[30][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[30][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[30][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[30][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[30][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[30][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[30][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[30][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[30][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[30][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[30][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[30][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[30][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[30][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[30][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[30][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[30][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[30][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[30][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[30][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[30][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[30][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[30][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[30][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[30][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[30][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[30][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[30][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[30][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[30][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[30][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[30][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[30][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[30][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[30][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[30][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[30][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[30][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[30][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[30][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[30][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[30][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[30][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[30][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[30][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[30][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[30][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[30][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[30][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[30][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[30][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[30][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[30][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[30][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[30][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[30][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[30][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[30][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[30][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[30][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[30][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[30][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[30][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[30][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[30][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[30][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[30][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 30, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[30][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[30][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[30][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[30][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[30][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[30].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[30][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[31][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[31][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[31][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[31][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[31][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[31][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[31][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[31][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[31][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[31][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[31][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[31][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[31][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[31][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[31][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[31][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[31][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[31][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[31][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[31][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[31][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[31][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[31][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[31][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[31][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[31][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[31][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[31][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[31][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[31][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[31][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[31][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[31][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[31][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[31][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[31][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[31][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[31][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[31][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[31][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[31][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[31][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[31][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[31][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[31][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[31][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[31][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[31][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[31][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[31][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[31][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[31][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[31][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[31][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[31][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[31][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[31][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[31][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[31][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[31][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[31][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[31][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[31][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[31][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[31][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[31][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[31][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[31][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[31][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[31][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[31][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[31][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[31][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[31][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[31][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[31][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[31][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[31][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[31][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[31][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[31][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[31][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[31][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[31][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[31][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[31][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[31][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[31][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[31][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[31][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[31][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[31][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[31][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[31][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[31][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[31][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[31][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[31][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[31][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[31][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[31][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[31][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[31][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[31][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[31][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[31][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[31][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[31][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[31][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[31][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[31][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[31][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[31][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[31][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[31][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[31][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[31][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[31][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[31][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[31][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[31][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[31][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[31][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[31][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[31][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[31][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[31][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[31][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[31][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[31][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[31][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[31][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[31][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[31][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[31][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[31][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[31][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[31][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[31][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[31][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[31][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[31][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[31][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[31][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[31][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[31][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[31][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[31][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[31][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[31][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[31][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[31][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[31][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[31][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[31][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[31][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[31][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[31][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[31][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[31][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[31][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[31][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[31][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[31][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[31][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[31][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[31][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[31][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[31][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[31][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[31][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[31][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[31][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[31][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[31][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[31][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[31][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[31][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[31][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[31][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[31][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[31][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[31][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[31][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[31][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[31][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 31, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[31][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[31][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[31][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[31][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[31][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[31].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[31][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[32][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[32][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[32][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[32][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[32][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[32][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[32][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[32][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[32][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[32][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[32][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[32][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[32][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[32][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[32][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[32][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[32][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[32][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[32][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[32][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[32][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[32][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[32][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[32][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[32][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[32][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[32][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[32][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[32][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[32][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[32][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[32][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[32][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[32][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[32][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[32][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[32][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[32][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[32][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[32][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[32][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[32][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[32][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[32][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[32][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[32][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[32][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[32][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[32][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[32][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[32][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[32][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[32][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[32][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[32][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[32][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[32][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[32][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[32][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[32][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[32][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[32][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[32][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[32][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[32][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[32][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[32][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[32][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[32][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[32][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[32][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[32][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[32][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[32][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[32][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[32][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[32][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[32][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[32][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[32][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[32][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[32][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[32][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[32][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[32][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[32][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[32][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[32][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[32][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[32][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[32][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[32][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[32][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[32][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[32][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[32][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[32][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[32][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[32][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[32][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[32][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[32][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[32][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[32][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[32][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[32][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[32][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[32][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[32][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[32][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[32][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[32][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[32][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[32][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[32][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[32][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[32][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[32][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[32][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[32][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[32][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[32][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[32][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[32][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[32][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[32][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[32][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[32][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[32][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[32][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[32][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[32][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[32][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[32][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[32][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[32][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[32][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[32][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[32][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[32][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[32][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[32][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[32][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[32][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[32][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[32][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[32][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[32][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[32][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[32][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[32][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[32][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[32][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[32][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[32][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[32][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[32][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[32][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[32][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[32][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[32][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[32][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[32][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[32][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[32][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[32][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[32][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[32][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[32][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[32][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[32][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[32][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[32][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[32][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[32][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[32][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[32][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[32][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[32][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[32][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[32][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[32][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[32][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[32][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[32][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[32][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 32, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[32][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[32][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[32][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[32][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[32][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[32].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[32][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[33][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[33][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[33][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[33][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[33][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[33][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[33][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[33][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[33][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[33][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[33][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[33][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[33][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[33][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[33][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[33][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[33][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[33][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[33][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[33][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[33][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[33][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[33][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[33][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[33][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[33][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[33][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[33][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[33][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[33][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[33][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[33][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[33][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[33][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[33][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[33][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[33][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[33][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[33][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[33][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[33][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[33][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[33][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[33][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[33][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[33][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[33][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[33][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[33][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[33][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[33][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[33][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[33][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[33][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[33][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[33][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[33][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[33][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[33][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[33][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[33][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[33][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[33][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[33][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[33][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[33][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[33][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[33][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[33][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[33][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[33][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[33][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[33][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[33][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[33][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[33][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[33][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[33][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[33][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[33][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[33][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[33][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[33][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[33][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[33][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[33][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[33][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[33][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[33][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[33][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[33][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[33][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[33][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[33][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[33][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[33][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[33][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[33][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[33][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[33][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[33][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[33][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[33][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[33][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[33][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[33][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[33][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[33][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[33][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[33][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[33][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[33][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[33][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[33][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[33][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[33][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[33][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[33][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[33][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[33][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[33][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[33][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[33][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[33][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[33][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[33][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[33][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[33][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[33][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[33][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[33][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[33][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[33][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[33][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[33][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[33][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[33][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[33][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[33][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[33][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[33][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[33][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[33][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[33][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[33][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[33][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[33][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[33][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[33][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[33][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[33][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[33][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[33][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[33][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[33][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[33][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[33][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[33][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[33][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[33][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[33][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[33][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[33][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[33][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[33][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[33][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[33][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[33][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[33][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[33][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[33][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[33][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[33][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[33][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[33][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[33][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[33][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[33][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[33][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[33][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[33][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[33][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[33][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[33][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[33][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[33][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 33, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[33][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[33][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[33][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[33][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[33][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[33].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[33][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[34][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[34][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[34][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[34][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[34][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[34][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[34][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[34][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[34][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[34][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[34][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[34][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[34][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[34][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[34][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[34][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[34][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[34][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[34][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[34][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[34][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[34][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[34][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[34][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[34][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[34][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[34][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[34][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[34][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[34][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[34][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[34][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[34][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[34][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[34][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[34][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[34][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[34][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[34][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[34][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[34][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[34][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[34][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[34][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[34][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[34][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[34][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[34][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[34][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[34][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[34][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[34][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[34][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[34][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[34][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[34][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[34][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[34][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[34][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[34][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[34][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[34][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[34][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[34][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[34][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[34][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[34][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[34][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[34][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[34][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[34][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[34][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[34][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[34][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[34][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[34][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[34][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[34][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[34][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[34][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[34][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[34][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[34][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[34][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[34][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[34][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[34][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[34][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[34][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[34][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[34][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[34][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[34][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[34][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[34][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[34][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[34][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[34][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[34][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[34][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[34][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[34][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[34][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[34][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[34][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[34][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[34][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[34][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[34][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[34][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[34][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[34][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[34][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[34][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[34][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[34][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[34][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[34][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[34][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[34][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[34][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[34][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[34][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[34][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[34][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[34][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[34][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[34][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[34][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[34][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[34][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[34][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[34][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[34][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[34][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[34][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[34][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[34][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[34][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[34][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[34][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[34][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[34][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[34][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[34][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[34][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[34][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[34][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[34][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[34][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[34][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[34][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[34][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[34][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[34][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[34][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[34][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[34][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[34][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[34][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[34][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[34][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[34][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[34][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[34][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[34][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[34][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[34][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[34][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[34][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[34][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[34][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[34][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[34][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[34][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[34][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[34][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[34][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[34][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[34][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[34][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[34][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[34][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[34][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[34][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[34][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 34, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[34][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[34][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[34][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[34][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[34][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[34].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[34][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[35][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[35][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[35][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[35][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[35][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[35][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[35][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[35][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[35][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[35][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[35][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[35][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[35][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[35][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[35][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[35][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[35][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[35][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[35][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[35][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[35][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[35][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[35][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[35][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[35][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[35][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[35][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[35][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[35][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[35][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[35][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[35][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[35][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[35][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[35][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[35][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[35][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[35][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[35][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[35][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[35][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[35][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[35][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[35][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[35][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[35][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[35][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[35][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[35][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[35][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[35][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[35][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[35][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[35][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[35][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[35][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[35][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[35][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[35][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[35][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[35][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[35][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[35][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[35][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[35][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[35][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[35][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[35][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[35][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[35][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[35][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[35][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[35][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[35][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[35][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[35][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[35][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[35][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[35][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[35][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[35][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[35][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[35][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[35][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[35][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[35][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[35][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[35][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[35][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[35][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[35][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[35][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[35][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[35][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[35][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[35][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[35][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[35][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[35][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[35][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[35][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[35][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[35][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[35][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[35][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[35][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[35][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[35][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[35][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[35][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[35][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[35][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[35][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[35][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[35][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[35][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[35][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[35][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[35][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[35][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[35][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[35][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[35][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[35][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[35][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[35][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[35][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[35][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[35][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[35][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[35][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[35][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[35][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[35][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[35][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[35][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[35][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[35][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[35][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[35][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[35][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[35][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[35][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[35][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[35][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[35][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[35][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[35][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[35][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[35][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[35][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[35][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[35][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[35][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[35][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[35][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[35][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[35][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[35][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[35][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[35][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[35][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[35][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[35][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[35][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[35][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[35][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[35][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[35][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[35][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[35][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[35][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[35][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[35][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[35][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[35][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[35][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[35][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[35][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[35][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[35][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[35][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[35][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[35][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[35][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[35][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 35, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[35][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[35][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[35][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[35][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[35][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[35].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[35][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[36][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[36][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[36][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[36][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[36][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[36][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[36][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[36][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[36][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[36][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[36][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[36][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[36][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[36][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[36][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[36][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[36][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[36][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[36][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[36][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[36][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[36][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[36][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[36][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[36][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[36][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[36][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[36][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[36][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[36][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[36][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[36][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[36][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[36][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[36][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[36][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[36][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[36][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[36][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[36][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[36][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[36][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[36][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[36][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[36][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[36][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[36][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[36][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[36][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[36][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[36][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[36][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[36][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[36][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[36][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[36][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[36][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[36][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[36][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[36][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[36][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[36][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[36][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[36][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[36][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[36][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[36][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[36][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[36][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[36][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[36][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[36][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[36][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[36][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[36][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[36][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[36][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[36][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[36][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[36][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[36][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[36][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[36][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[36][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[36][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[36][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[36][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[36][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[36][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[36][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[36][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[36][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[36][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[36][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[36][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[36][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[36][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[36][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[36][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[36][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[36][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[36][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[36][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[36][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[36][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[36][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[36][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[36][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[36][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[36][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[36][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[36][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[36][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[36][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[36][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[36][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[36][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[36][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[36][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[36][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[36][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[36][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[36][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[36][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[36][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[36][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[36][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[36][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[36][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[36][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[36][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[36][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[36][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[36][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[36][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[36][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[36][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[36][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[36][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[36][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[36][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[36][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[36][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[36][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[36][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[36][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[36][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[36][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[36][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[36][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[36][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[36][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[36][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[36][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[36][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[36][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[36][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[36][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[36][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[36][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[36][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[36][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[36][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[36][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[36][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[36][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[36][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[36][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[36][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[36][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[36][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[36][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[36][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[36][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[36][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[36][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[36][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[36][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[36][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[36][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[36][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[36][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[36][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[36][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[36][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[36][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 36, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[36][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[36][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[36][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[36][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[36][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[36].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[36][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[37][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[37][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[37][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[37][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[37][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[37][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[37][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[37][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[37][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[37][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[37][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[37][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[37][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[37][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[37][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[37][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[37][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[37][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[37][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[37][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[37][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[37][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[37][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[37][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[37][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[37][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[37][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[37][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[37][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[37][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[37][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[37][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[37][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[37][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[37][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[37][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[37][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[37][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[37][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[37][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[37][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[37][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[37][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[37][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[37][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[37][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[37][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[37][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[37][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[37][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[37][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[37][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[37][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[37][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[37][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[37][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[37][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[37][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[37][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[37][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[37][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[37][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[37][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[37][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[37][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[37][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[37][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[37][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[37][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[37][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[37][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[37][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[37][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[37][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[37][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[37][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[37][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[37][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[37][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[37][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[37][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[37][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[37][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[37][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[37][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[37][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[37][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[37][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[37][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[37][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[37][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[37][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[37][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[37][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[37][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[37][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[37][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[37][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[37][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[37][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[37][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[37][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[37][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[37][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[37][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[37][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[37][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[37][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[37][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[37][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[37][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[37][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[37][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[37][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[37][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[37][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[37][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[37][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[37][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[37][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[37][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[37][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[37][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[37][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[37][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[37][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[37][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[37][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[37][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[37][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[37][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[37][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[37][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[37][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[37][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[37][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[37][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[37][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[37][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[37][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[37][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[37][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[37][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[37][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[37][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[37][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[37][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[37][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[37][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[37][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[37][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[37][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[37][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[37][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[37][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[37][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[37][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[37][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[37][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[37][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[37][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[37][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[37][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[37][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[37][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[37][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[37][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[37][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[37][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[37][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[37][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[37][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[37][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[37][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[37][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[37][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[37][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[37][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[37][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[37][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[37][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[37][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[37][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[37][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[37][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[37][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 37, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[37][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[37][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[37][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[37][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[37][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[37].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[37][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[38][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[38][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[38][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[38][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[38][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[38][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[38][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[38][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[38][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[38][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[38][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[38][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[38][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[38][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[38][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[38][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[38][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[38][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[38][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[38][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[38][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[38][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[38][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[38][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[38][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[38][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[38][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[38][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[38][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[38][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[38][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[38][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[38][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[38][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[38][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[38][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[38][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[38][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[38][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[38][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[38][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[38][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[38][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[38][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[38][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[38][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[38][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[38][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[38][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[38][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[38][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[38][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[38][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[38][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[38][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[38][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[38][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[38][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[38][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[38][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[38][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[38][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[38][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[38][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[38][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[38][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[38][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[38][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[38][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[38][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[38][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[38][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[38][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[38][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[38][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[38][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[38][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[38][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[38][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[38][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[38][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[38][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[38][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[38][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[38][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[38][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[38][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[38][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[38][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[38][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[38][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[38][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[38][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[38][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[38][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[38][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[38][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[38][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[38][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[38][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[38][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[38][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[38][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[38][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[38][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[38][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[38][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[38][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[38][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[38][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[38][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[38][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[38][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[38][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[38][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[38][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[38][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[38][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[38][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[38][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[38][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[38][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[38][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[38][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[38][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[38][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[38][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[38][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[38][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[38][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[38][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[38][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[38][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[38][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[38][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[38][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[38][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[38][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[38][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[38][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[38][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[38][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[38][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[38][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[38][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[38][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[38][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[38][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[38][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[38][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[38][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[38][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[38][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[38][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[38][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[38][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[38][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[38][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[38][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[38][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[38][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[38][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[38][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[38][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[38][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[38][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[38][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[38][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[38][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[38][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[38][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[38][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[38][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[38][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[38][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[38][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[38][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[38][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[38][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[38][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[38][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[38][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[38][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[38][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[38][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[38][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 38, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[38][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[38][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[38][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[38][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[38][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[38].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[38][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[39][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[39][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[39][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[39][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[39][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[39][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[39][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[39][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[39][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[39][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[39][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[39][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[39][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[39][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[39][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[39][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[39][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[39][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[39][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[39][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[39][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[39][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[39][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[39][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[39][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[39][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[39][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[39][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[39][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[39][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[39][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[39][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[39][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[39][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[39][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[39][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[39][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[39][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[39][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[39][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[39][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[39][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[39][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[39][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[39][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[39][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[39][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[39][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[39][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[39][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[39][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[39][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[39][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[39][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[39][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[39][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[39][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[39][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[39][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[39][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[39][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[39][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[39][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[39][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[39][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[39][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[39][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[39][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[39][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[39][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[39][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[39][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[39][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[39][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[39][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[39][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[39][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[39][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[39][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[39][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[39][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[39][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[39][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[39][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[39][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[39][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[39][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[39][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[39][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[39][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[39][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[39][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[39][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[39][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[39][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[39][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[39][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[39][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[39][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[39][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[39][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[39][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[39][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[39][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[39][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[39][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[39][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[39][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[39][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[39][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[39][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[39][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[39][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[39][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[39][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[39][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[39][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[39][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[39][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[39][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[39][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[39][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[39][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[39][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[39][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[39][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[39][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[39][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[39][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[39][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[39][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[39][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[39][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[39][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[39][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[39][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[39][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[39][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[39][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[39][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[39][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[39][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[39][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[39][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[39][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[39][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[39][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[39][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[39][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[39][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[39][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[39][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[39][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[39][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[39][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[39][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[39][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[39][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[39][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[39][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[39][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[39][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[39][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[39][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[39][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[39][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[39][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[39][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[39][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[39][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[39][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[39][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[39][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[39][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[39][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[39][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[39][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[39][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[39][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[39][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[39][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[39][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[39][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[39][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[39][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[39][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 39, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[39][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[39][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[39][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[39][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[39][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[39].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[39][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[40][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[40][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[40][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[40][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[40][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[40][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[40][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[40][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[40][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[40][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[40][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[40][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[40][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[40][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[40][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[40][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[40][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[40][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[40][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[40][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[40][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[40][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[40][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[40][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[40][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[40][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[40][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[40][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[40][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[40][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[40][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[40][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[40][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[40][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[40][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[40][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[40][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[40][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[40][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[40][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[40][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[40][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[40][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[40][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[40][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[40][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[40][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[40][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[40][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[40][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[40][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[40][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[40][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[40][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[40][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[40][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[40][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[40][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[40][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[40][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[40][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[40][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[40][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[40][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[40][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[40][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[40][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[40][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[40][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[40][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[40][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[40][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[40][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[40][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[40][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[40][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[40][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[40][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[40][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[40][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[40][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[40][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[40][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[40][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[40][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[40][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[40][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[40][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[40][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[40][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[40][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[40][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[40][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[40][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[40][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[40][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[40][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[40][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[40][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[40][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[40][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[40][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[40][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[40][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[40][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[40][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[40][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[40][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[40][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[40][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[40][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[40][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[40][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[40][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[40][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[40][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[40][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[40][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[40][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[40][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[40][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[40][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[40][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[40][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[40][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[40][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[40][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[40][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[40][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[40][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[40][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[40][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[40][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[40][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[40][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[40][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[40][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[40][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[40][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[40][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[40][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[40][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[40][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[40][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[40][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[40][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[40][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[40][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[40][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[40][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[40][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[40][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[40][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[40][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[40][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[40][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[40][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[40][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[40][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[40][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[40][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[40][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[40][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[40][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[40][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[40][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[40][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[40][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[40][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[40][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[40][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[40][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[40][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[40][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[40][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[40][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[40][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[40][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[40][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[40][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[40][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[40][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[40][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[40][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[40][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[40][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 40, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[40][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[40][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[40][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[40][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[40][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[40].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[40][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[41][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[41][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[41][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[41][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[41][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[41][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[41][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[41][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[41][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[41][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[41][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[41][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[41][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[41][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[41][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[41][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[41][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[41][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[41][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[41][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[41][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[41][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[41][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[41][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[41][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[41][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[41][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[41][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[41][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[41][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[41][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[41][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[41][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[41][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[41][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[41][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[41][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[41][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[41][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[41][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[41][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[41][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[41][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[41][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[41][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[41][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[41][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[41][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[41][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[41][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[41][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[41][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[41][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[41][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[41][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[41][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[41][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[41][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[41][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[41][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[41][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[41][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[41][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[41][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[41][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[41][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[41][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[41][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[41][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[41][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[41][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[41][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[41][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[41][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[41][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[41][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[41][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[41][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[41][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[41][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[41][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[41][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[41][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[41][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[41][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[41][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[41][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[41][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[41][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[41][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[41][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[41][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[41][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[41][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[41][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[41][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[41][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[41][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[41][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[41][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[41][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[41][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[41][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[41][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[41][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[41][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[41][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[41][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[41][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[41][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[41][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[41][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[41][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[41][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[41][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[41][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[41][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[41][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[41][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[41][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[41][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[41][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[41][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[41][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[41][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[41][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[41][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[41][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[41][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[41][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[41][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[41][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[41][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[41][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[41][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[41][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[41][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[41][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[41][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[41][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[41][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[41][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[41][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[41][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[41][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[41][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[41][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[41][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[41][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[41][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[41][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[41][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[41][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[41][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[41][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[41][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[41][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[41][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[41][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[41][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[41][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[41][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[41][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[41][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[41][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[41][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[41][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[41][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[41][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[41][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[41][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[41][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[41][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[41][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[41][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[41][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[41][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[41][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[41][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[41][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[41][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[41][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[41][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[41][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[41][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[41][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 41, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[41][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[41][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[41][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[41][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[41][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[41].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[41][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[42][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[42][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[42][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[42][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[42][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[42][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[42][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[42][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[42][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[42][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[42][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[42][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[42][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[42][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[42][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[42][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[42][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[42][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[42][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[42][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[42][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[42][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[42][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[42][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[42][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[42][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[42][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[42][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[42][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[42][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[42][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[42][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[42][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[42][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[42][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[42][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[42][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[42][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[42][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[42][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[42][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[42][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[42][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[42][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[42][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[42][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[42][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[42][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[42][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[42][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[42][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[42][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[42][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[42][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[42][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[42][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[42][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[42][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[42][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[42][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[42][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[42][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[42][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[42][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[42][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[42][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[42][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[42][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[42][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[42][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[42][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[42][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[42][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[42][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[42][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[42][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[42][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[42][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[42][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[42][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[42][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[42][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[42][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[42][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[42][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[42][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[42][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[42][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[42][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[42][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[42][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[42][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[42][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[42][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[42][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[42][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[42][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[42][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[42][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[42][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[42][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[42][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[42][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[42][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[42][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[42][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[42][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[42][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[42][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[42][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[42][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[42][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[42][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[42][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[42][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[42][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[42][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[42][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[42][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[42][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[42][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[42][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[42][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[42][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[42][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[42][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[42][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[42][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[42][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[42][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[42][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[42][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[42][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[42][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[42][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[42][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[42][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[42][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[42][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[42][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[42][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[42][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[42][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[42][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[42][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[42][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[42][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[42][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[42][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[42][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[42][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[42][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[42][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[42][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[42][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[42][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[42][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[42][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[42][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[42][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[42][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[42][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[42][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[42][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[42][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[42][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[42][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[42][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[42][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[42][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[42][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[42][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[42][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[42][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[42][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[42][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[42][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[42][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[42][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[42][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[42][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[42][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[42][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[42][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[42][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[42][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 42, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[42][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[42][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[42][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[42][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[42][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[42].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[42][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[43][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[43][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[43][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[43][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[43][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[43][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[43][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[43][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[43][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[43][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[43][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[43][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[43][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[43][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[43][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[43][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[43][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[43][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[43][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[43][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[43][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[43][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[43][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[43][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[43][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[43][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[43][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[43][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[43][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[43][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[43][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[43][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[43][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[43][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[43][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[43][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[43][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[43][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[43][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[43][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[43][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[43][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[43][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[43][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[43][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[43][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[43][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[43][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[43][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[43][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[43][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[43][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[43][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[43][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[43][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[43][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[43][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[43][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[43][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[43][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[43][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[43][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[43][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[43][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[43][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[43][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[43][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[43][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[43][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[43][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[43][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[43][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[43][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[43][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[43][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[43][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[43][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[43][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[43][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[43][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[43][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[43][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[43][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[43][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[43][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[43][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[43][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[43][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[43][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[43][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[43][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[43][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[43][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[43][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[43][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[43][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[43][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[43][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[43][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[43][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[43][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[43][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[43][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[43][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[43][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[43][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[43][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[43][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[43][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[43][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[43][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[43][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[43][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[43][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[43][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[43][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[43][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[43][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[43][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[43][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[43][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[43][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[43][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[43][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[43][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[43][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[43][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[43][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[43][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[43][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[43][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[43][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[43][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[43][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[43][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[43][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[43][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[43][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[43][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[43][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[43][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[43][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[43][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[43][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[43][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[43][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[43][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[43][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[43][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[43][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[43][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[43][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[43][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[43][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[43][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[43][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[43][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[43][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[43][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[43][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[43][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[43][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[43][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[43][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[43][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[43][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[43][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[43][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[43][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[43][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[43][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[43][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[43][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[43][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[43][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[43][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[43][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[43][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[43][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[43][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[43][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[43][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[43][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[43][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[43][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[43][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 43, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[43][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[43][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[43][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[43][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[43][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[43].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[43][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[44][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[44][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[44][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[44][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[44][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[44][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[44][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[44][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[44][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[44][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[44][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[44][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[44][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[44][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[44][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[44][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[44][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[44][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[44][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[44][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[44][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[44][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[44][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[44][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[44][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[44][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[44][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[44][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[44][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[44][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[44][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[44][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[44][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[44][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[44][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[44][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[44][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[44][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[44][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[44][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[44][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[44][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[44][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[44][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[44][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[44][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[44][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[44][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[44][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[44][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[44][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[44][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[44][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[44][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[44][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[44][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[44][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[44][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[44][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[44][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[44][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[44][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[44][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[44][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[44][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[44][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[44][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[44][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[44][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[44][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[44][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[44][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[44][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[44][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[44][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[44][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[44][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[44][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[44][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[44][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[44][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[44][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[44][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[44][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[44][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[44][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[44][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[44][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[44][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[44][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[44][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[44][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[44][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[44][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[44][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[44][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[44][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[44][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[44][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[44][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[44][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[44][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[44][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[44][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[44][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[44][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[44][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[44][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[44][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[44][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[44][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[44][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[44][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[44][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[44][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[44][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[44][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[44][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[44][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[44][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[44][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[44][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[44][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[44][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[44][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[44][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[44][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[44][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[44][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[44][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[44][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[44][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[44][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[44][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[44][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[44][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[44][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[44][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[44][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[44][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[44][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[44][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[44][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[44][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[44][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[44][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[44][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[44][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[44][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[44][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[44][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[44][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[44][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[44][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[44][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[44][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[44][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[44][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[44][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[44][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[44][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[44][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[44][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[44][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[44][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[44][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[44][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[44][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[44][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[44][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[44][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[44][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[44][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[44][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[44][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[44][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[44][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[44][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[44][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[44][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[44][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[44][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[44][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[44][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[44][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[44][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 44, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[44][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[44][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[44][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[44][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[44][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[44].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[44][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[45][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[45][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[45][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[45][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[45][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[45][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[45][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[45][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[45][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[45][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[45][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[45][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[45][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[45][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[45][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[45][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[45][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[45][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[45][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[45][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[45][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[45][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[45][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[45][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[45][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[45][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[45][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[45][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[45][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[45][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[45][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[45][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[45][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[45][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[45][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[45][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[45][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[45][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[45][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[45][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[45][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[45][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[45][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[45][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[45][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[45][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[45][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[45][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[45][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[45][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[45][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[45][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[45][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[45][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[45][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[45][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[45][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[45][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[45][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[45][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[45][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[45][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[45][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[45][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[45][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[45][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[45][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[45][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[45][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[45][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[45][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[45][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[45][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[45][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[45][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[45][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[45][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[45][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[45][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[45][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[45][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[45][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[45][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[45][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[45][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[45][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[45][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[45][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[45][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[45][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[45][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[45][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[45][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[45][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[45][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[45][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[45][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[45][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[45][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[45][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[45][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[45][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[45][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[45][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[45][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[45][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[45][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[45][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[45][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[45][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[45][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[45][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[45][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[45][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[45][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[45][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[45][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[45][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[45][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[45][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[45][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[45][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[45][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[45][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[45][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[45][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[45][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[45][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[45][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[45][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[45][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[45][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[45][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[45][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[45][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[45][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[45][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[45][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[45][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[45][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[45][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[45][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[45][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[45][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[45][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[45][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[45][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[45][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[45][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[45][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[45][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[45][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[45][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[45][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[45][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[45][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[45][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[45][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[45][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[45][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[45][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[45][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[45][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[45][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[45][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[45][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[45][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[45][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[45][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[45][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[45][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[45][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[45][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[45][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[45][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[45][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[45][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[45][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[45][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[45][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[45][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[45][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[45][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[45][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[45][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[45][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 45, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[45][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[45][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[45][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[45][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[45][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[45].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[45][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[46][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[46][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[46][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[46][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[46][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[46][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[46][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[46][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[46][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[46][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[46][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[46][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[46][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[46][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[46][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[46][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[46][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[46][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[46][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[46][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[46][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[46][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[46][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[46][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[46][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[46][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[46][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[46][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[46][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[46][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[46][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[46][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[46][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[46][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[46][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[46][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[46][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[46][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[46][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[46][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[46][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[46][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[46][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[46][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[46][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[46][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[46][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[46][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[46][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[46][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[46][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[46][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[46][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[46][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[46][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[46][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[46][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[46][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[46][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[46][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[46][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[46][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[46][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[46][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[46][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[46][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[46][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[46][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[46][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[46][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[46][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[46][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[46][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[46][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[46][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[46][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[46][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[46][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[46][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[46][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[46][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[46][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[46][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[46][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[46][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[46][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[46][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[46][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[46][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[46][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[46][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[46][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[46][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[46][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[46][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[46][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[46][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[46][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[46][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[46][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[46][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[46][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[46][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[46][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[46][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[46][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[46][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[46][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[46][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[46][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[46][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[46][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[46][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[46][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[46][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[46][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[46][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[46][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[46][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[46][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[46][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[46][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[46][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[46][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[46][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[46][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[46][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[46][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[46][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[46][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[46][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[46][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[46][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[46][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[46][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[46][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[46][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[46][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[46][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[46][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[46][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[46][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[46][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[46][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[46][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[46][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[46][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[46][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[46][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[46][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[46][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[46][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[46][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[46][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[46][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[46][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[46][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[46][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[46][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[46][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[46][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[46][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[46][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[46][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[46][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[46][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[46][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[46][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[46][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[46][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[46][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[46][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[46][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[46][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[46][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[46][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[46][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[46][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[46][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[46][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[46][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[46][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[46][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[46][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[46][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[46][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 46, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[46][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[46][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[46][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[46][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[46][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[46].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[46][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[47][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[47][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[47][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[47][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[47][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[47][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[47][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[47][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[47][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[47][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[47][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[47][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[47][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[47][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[47][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[47][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[47][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[47][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[47][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[47][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[47][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[47][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[47][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[47][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[47][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[47][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[47][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[47][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[47][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[47][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[47][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[47][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[47][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[47][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[47][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[47][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[47][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[47][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[47][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[47][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[47][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[47][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[47][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[47][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[47][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[47][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[47][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[47][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[47][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[47][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[47][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[47][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[47][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[47][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[47][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[47][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[47][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[47][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[47][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[47][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[47][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[47][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[47][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[47][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[47][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[47][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[47][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[47][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[47][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[47][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[47][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[47][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[47][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[47][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[47][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[47][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[47][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[47][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[47][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[47][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[47][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[47][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[47][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[47][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[47][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[47][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[47][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[47][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[47][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[47][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[47][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[47][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[47][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[47][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[47][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[47][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[47][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[47][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[47][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[47][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[47][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[47][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[47][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[47][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[47][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[47][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[47][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[47][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[47][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[47][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[47][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[47][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[47][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[47][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[47][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[47][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[47][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[47][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[47][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[47][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[47][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[47][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[47][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[47][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[47][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[47][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[47][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[47][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[47][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[47][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[47][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[47][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[47][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[47][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[47][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[47][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[47][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[47][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[47][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[47][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[47][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[47][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[47][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[47][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[47][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[47][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[47][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[47][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[47][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[47][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[47][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[47][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[47][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[47][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[47][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[47][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[47][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[47][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[47][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[47][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[47][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[47][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[47][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[47][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[47][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[47][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[47][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[47][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[47][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[47][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[47][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[47][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[47][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[47][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[47][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[47][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[47][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[47][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[47][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[47][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[47][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[47][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[47][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[47][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[47][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[47][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 47, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[47][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[47][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[47][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[47][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[47][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[47].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[47][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[48][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[48][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[48][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[48][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[48][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[48][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[48][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[48][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[48][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[48][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[48][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[48][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[48][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[48][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[48][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[48][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[48][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[48][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[48][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[48][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[48][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[48][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[48][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[48][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[48][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[48][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[48][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[48][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[48][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[48][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[48][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[48][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[48][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[48][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[48][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[48][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[48][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[48][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[48][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[48][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[48][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[48][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[48][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[48][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[48][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[48][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[48][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[48][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[48][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[48][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[48][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[48][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[48][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[48][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[48][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[48][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[48][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[48][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[48][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[48][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[48][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[48][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[48][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[48][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[48][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[48][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[48][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[48][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[48][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[48][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[48][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[48][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[48][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[48][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[48][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[48][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[48][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[48][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[48][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[48][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[48][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[48][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[48][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[48][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[48][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[48][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[48][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[48][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[48][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[48][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[48][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[48][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[48][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[48][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[48][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[48][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[48][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[48][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[48][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[48][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[48][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[48][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[48][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[48][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[48][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[48][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[48][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[48][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[48][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[48][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[48][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[48][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[48][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[48][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[48][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[48][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[48][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[48][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[48][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[48][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[48][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[48][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[48][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[48][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[48][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[48][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[48][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[48][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[48][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[48][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[48][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[48][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[48][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[48][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[48][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[48][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[48][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[48][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[48][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[48][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[48][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[48][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[48][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[48][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[48][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[48][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[48][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[48][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[48][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[48][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[48][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[48][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[48][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[48][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[48][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[48][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[48][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[48][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[48][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[48][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[48][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[48][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[48][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[48][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[48][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[48][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[48][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[48][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[48][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[48][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[48][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[48][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[48][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[48][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[48][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[48][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[48][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[48][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[48][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[48][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[48][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[48][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[48][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[48][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[48][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[48][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 48, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[48][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[48][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[48][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[48][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[48][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[48].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[48][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[49][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[49][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[49][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[49][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[49][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[49][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[49][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[49][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[49][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[49][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[49][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[49][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[49][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[49][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[49][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[49][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[49][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[49][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[49][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[49][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[49][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[49][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[49][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[49][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[49][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[49][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[49][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[49][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[49][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[49][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[49][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[49][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[49][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[49][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[49][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[49][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[49][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[49][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[49][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[49][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[49][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[49][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[49][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[49][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[49][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[49][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[49][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[49][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[49][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[49][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[49][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[49][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[49][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[49][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[49][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[49][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[49][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[49][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[49][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[49][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[49][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[49][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[49][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[49][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[49][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[49][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[49][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[49][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[49][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[49][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[49][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[49][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[49][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[49][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[49][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[49][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[49][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[49][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[49][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[49][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[49][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[49][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[49][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[49][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[49][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[49][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[49][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[49][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[49][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[49][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[49][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[49][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[49][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[49][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[49][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[49][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[49][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[49][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[49][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[49][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[49][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[49][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[49][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[49][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[49][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[49][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[49][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[49][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[49][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[49][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[49][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[49][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[49][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[49][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[49][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[49][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[49][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[49][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[49][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[49][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[49][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[49][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[49][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[49][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[49][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[49][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[49][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[49][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[49][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[49][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[49][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[49][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[49][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[49][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[49][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[49][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[49][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[49][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[49][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[49][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[49][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[49][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[49][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[49][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[49][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[49][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[49][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[49][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[49][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[49][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[49][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[49][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[49][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[49][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[49][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[49][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[49][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[49][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[49][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[49][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[49][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[49][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[49][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[49][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[49][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[49][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[49][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[49][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[49][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[49][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[49][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[49][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[49][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[49][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[49][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[49][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[49][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[49][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[49][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[49][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[49][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[49][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[49][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[49][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[49][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[49][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 49, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[49][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[49][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[49][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[49][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[49][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[49].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[49][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[50][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[50][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[50][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[50][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[50][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[50][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[50][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[50][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[50][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[50][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[50][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[50][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[50][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[50][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[50][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[50][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[50][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[50][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[50][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[50][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[50][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[50][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[50][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[50][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[50][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[50][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[50][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[50][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[50][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[50][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[50][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[50][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[50][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[50][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[50][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[50][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[50][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[50][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[50][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[50][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[50][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[50][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[50][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[50][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[50][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[50][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[50][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[50][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[50][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[50][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[50][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[50][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[50][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[50][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[50][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[50][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[50][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[50][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[50][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[50][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[50][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[50][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[50][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[50][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[50][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[50][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[50][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[50][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[50][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[50][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[50][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[50][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[50][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[50][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[50][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[50][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[50][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[50][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[50][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[50][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[50][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[50][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[50][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[50][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[50][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[50][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[50][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[50][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[50][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[50][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[50][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[50][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[50][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[50][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[50][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[50][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[50][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[50][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[50][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[50][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[50][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[50][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[50][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[50][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[50][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[50][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[50][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[50][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[50][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[50][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[50][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[50][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[50][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[50][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[50][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[50][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[50][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[50][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[50][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[50][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[50][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[50][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[50][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[50][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[50][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[50][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[50][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[50][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[50][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[50][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[50][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[50][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[50][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[50][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[50][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[50][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[50][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[50][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[50][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[50][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[50][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[50][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[50][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[50][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[50][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[50][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[50][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[50][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[50][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[50][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[50][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[50][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[50][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[50][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[50][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[50][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[50][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[50][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[50][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[50][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[50][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[50][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[50][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[50][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[50][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[50][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[50][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[50][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[50][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[50][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[50][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[50][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[50][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[50][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[50][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[50][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[50][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[50][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[50][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[50][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[50][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[50][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[50][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[50][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[50][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[50][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 50, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[50][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[50][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[50][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[50][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[50][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[50].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[50][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[51][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[51][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[51][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[51][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[51][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[51][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[51][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[51][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[51][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[51][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[51][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[51][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[51][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[51][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[51][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[51][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[51][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[51][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[51][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[51][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[51][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[51][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[51][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[51][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[51][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[51][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[51][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[51][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[51][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[51][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[51][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[51][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[51][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[51][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[51][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[51][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[51][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[51][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[51][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[51][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[51][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[51][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[51][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[51][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[51][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[51][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[51][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[51][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[51][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[51][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[51][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[51][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[51][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[51][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[51][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[51][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[51][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[51][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[51][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[51][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[51][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[51][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[51][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[51][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[51][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[51][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[51][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[51][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[51][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[51][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[51][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[51][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[51][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[51][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[51][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[51][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[51][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[51][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[51][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[51][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[51][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[51][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[51][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[51][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[51][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[51][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[51][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[51][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[51][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[51][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[51][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[51][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[51][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[51][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[51][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[51][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[51][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[51][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[51][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[51][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[51][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[51][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[51][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[51][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[51][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[51][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[51][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[51][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[51][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[51][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[51][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[51][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[51][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[51][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[51][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[51][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[51][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[51][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[51][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[51][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[51][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[51][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[51][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[51][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[51][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[51][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[51][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[51][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[51][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[51][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[51][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[51][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[51][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[51][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[51][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[51][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[51][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[51][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[51][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[51][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[51][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[51][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[51][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[51][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[51][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[51][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[51][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[51][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[51][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[51][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[51][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[51][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[51][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[51][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[51][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[51][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[51][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[51][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[51][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[51][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[51][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[51][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[51][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[51][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[51][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[51][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[51][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[51][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[51][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[51][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[51][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[51][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[51][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[51][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[51][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[51][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[51][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[51][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[51][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[51][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[51][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[51][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[51][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[51][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[51][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[51][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 51, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[51][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[51][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[51][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[51][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[51][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[51].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[51][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[52][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[52][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[52][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[52][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[52][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[52][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[52][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[52][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[52][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[52][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[52][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[52][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[52][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[52][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[52][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[52][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[52][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[52][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[52][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[52][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[52][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[52][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[52][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[52][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[52][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[52][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[52][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[52][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[52][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[52][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[52][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[52][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[52][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[52][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[52][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[52][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[52][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[52][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[52][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[52][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[52][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[52][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[52][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[52][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[52][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[52][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[52][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[52][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[52][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[52][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[52][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[52][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[52][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[52][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[52][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[52][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[52][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[52][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[52][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[52][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[52][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[52][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[52][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[52][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[52][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[52][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[52][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[52][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[52][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[52][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[52][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[52][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[52][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[52][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[52][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[52][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[52][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[52][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[52][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[52][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[52][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[52][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[52][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[52][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[52][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[52][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[52][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[52][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[52][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[52][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[52][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[52][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[52][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[52][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[52][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[52][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[52][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[52][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[52][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[52][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[52][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[52][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[52][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[52][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[52][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[52][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[52][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[52][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[52][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[52][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[52][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[52][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[52][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[52][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[52][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[52][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[52][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[52][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[52][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[52][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[52][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[52][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[52][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[52][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[52][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[52][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[52][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[52][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[52][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[52][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[52][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[52][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[52][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[52][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[52][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[52][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[52][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[52][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[52][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[52][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[52][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[52][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[52][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[52][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[52][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[52][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[52][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[52][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[52][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[52][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[52][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[52][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[52][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[52][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[52][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[52][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[52][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[52][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[52][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[52][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[52][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[52][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[52][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[52][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[52][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[52][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[52][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[52][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[52][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[52][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[52][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[52][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[52][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[52][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[52][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[52][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[52][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[52][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[52][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[52][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[52][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[52][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[52][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[52][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[52][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[52][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 52, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[52][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[52][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[52][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[52][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[52][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[52].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[52][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[53][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[53][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[53][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[53][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[53][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[53][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[53][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[53][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[53][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[53][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[53][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[53][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[53][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[53][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[53][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[53][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[53][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[53][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[53][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[53][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[53][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[53][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[53][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[53][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[53][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[53][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[53][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[53][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[53][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[53][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[53][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[53][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[53][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[53][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[53][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[53][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[53][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[53][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[53][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[53][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[53][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[53][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[53][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[53][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[53][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[53][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[53][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[53][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[53][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[53][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[53][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[53][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[53][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[53][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[53][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[53][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[53][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[53][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[53][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[53][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[53][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[53][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[53][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[53][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[53][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[53][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[53][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[53][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[53][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[53][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[53][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[53][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[53][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[53][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[53][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[53][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[53][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[53][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[53][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[53][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[53][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[53][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[53][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[53][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[53][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[53][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[53][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[53][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[53][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[53][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[53][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[53][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[53][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[53][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[53][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[53][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[53][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[53][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[53][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[53][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[53][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[53][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[53][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[53][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[53][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[53][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[53][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[53][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[53][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[53][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[53][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[53][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[53][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[53][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[53][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[53][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[53][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[53][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[53][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[53][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[53][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[53][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[53][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[53][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[53][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[53][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[53][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[53][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[53][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[53][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[53][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[53][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[53][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[53][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[53][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[53][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[53][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[53][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[53][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[53][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[53][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[53][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[53][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[53][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[53][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[53][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[53][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[53][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[53][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[53][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[53][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[53][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[53][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[53][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[53][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[53][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[53][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[53][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[53][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[53][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[53][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[53][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[53][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[53][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[53][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[53][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[53][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[53][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[53][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[53][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[53][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[53][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[53][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[53][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[53][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[53][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[53][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[53][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[53][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[53][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[53][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[53][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[53][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[53][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[53][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[53][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 53, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[53][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[53][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[53][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[53][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[53][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[53].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[53][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[54][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[54][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[54][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[54][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[54][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[54][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[54][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[54][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[54][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[54][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[54][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[54][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[54][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[54][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[54][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[54][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[54][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[54][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[54][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[54][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[54][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[54][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[54][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[54][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[54][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[54][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[54][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[54][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[54][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[54][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[54][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[54][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[54][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[54][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[54][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[54][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[54][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[54][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[54][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[54][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[54][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[54][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[54][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[54][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[54][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[54][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[54][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[54][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[54][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[54][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[54][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[54][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[54][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[54][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[54][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[54][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[54][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[54][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[54][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[54][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[54][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[54][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[54][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[54][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[54][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[54][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[54][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[54][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[54][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[54][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[54][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[54][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[54][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[54][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[54][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[54][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[54][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[54][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[54][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[54][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[54][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[54][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[54][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[54][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[54][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[54][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[54][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[54][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[54][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[54][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[54][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[54][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[54][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[54][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[54][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[54][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[54][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[54][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[54][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[54][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[54][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[54][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[54][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[54][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[54][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[54][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[54][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[54][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[54][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[54][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[54][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[54][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[54][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[54][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[54][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[54][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[54][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[54][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[54][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[54][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[54][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[54][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[54][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[54][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[54][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[54][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[54][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[54][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[54][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[54][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[54][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[54][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[54][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[54][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[54][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[54][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[54][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[54][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[54][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[54][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[54][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[54][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[54][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[54][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[54][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[54][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[54][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[54][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[54][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[54][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[54][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[54][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[54][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[54][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[54][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[54][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[54][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[54][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[54][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[54][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[54][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[54][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[54][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[54][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[54][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[54][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[54][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[54][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[54][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[54][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[54][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[54][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[54][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[54][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[54][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[54][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[54][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[54][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[54][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[54][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[54][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[54][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[54][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[54][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[54][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[54][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 54, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[54][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[54][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[54][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[54][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[54][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[54].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[54][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[55][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[55][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[55][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[55][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[55][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[55][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[55][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[55][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[55][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[55][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[55][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[55][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[55][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[55][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[55][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[55][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[55][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[55][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[55][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[55][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[55][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[55][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[55][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[55][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[55][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[55][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[55][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[55][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[55][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[55][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[55][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[55][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[55][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[55][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[55][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[55][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[55][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[55][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[55][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[55][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[55][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[55][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[55][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[55][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[55][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[55][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[55][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[55][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[55][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[55][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[55][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[55][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[55][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[55][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[55][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[55][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[55][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[55][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[55][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[55][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[55][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[55][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[55][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[55][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[55][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[55][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[55][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[55][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[55][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[55][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[55][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[55][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[55][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[55][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[55][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[55][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[55][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[55][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[55][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[55][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[55][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[55][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[55][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[55][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[55][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[55][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[55][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[55][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[55][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[55][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[55][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[55][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[55][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[55][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[55][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[55][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[55][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[55][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[55][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[55][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[55][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[55][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[55][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[55][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[55][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[55][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[55][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[55][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[55][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[55][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[55][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[55][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[55][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[55][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[55][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[55][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[55][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[55][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[55][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[55][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[55][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[55][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[55][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[55][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[55][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[55][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[55][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[55][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[55][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[55][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[55][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[55][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[55][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[55][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[55][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[55][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[55][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[55][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[55][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[55][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[55][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[55][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[55][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[55][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[55][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[55][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[55][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[55][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[55][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[55][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[55][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[55][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[55][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[55][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[55][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[55][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[55][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[55][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[55][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[55][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[55][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[55][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[55][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[55][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[55][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[55][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[55][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[55][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[55][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[55][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[55][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[55][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[55][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[55][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[55][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[55][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[55][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[55][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[55][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[55][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[55][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[55][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[55][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[55][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[55][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[55][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 55, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[55][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[55][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[55][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[55][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[55][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[55].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[55][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[56][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[56][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[56][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[56][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[56][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[56][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[56][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[56][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[56][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[56][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[56][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[56][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[56][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[56][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[56][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[56][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[56][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[56][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[56][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[56][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[56][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[56][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[56][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[56][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[56][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[56][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[56][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[56][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[56][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[56][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[56][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[56][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[56][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[56][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[56][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[56][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[56][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[56][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[56][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[56][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[56][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[56][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[56][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[56][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[56][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[56][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[56][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[56][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[56][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[56][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[56][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[56][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[56][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[56][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[56][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[56][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[56][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[56][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[56][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[56][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[56][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[56][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[56][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[56][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[56][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[56][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[56][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[56][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[56][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[56][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[56][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[56][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[56][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[56][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[56][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[56][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[56][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[56][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[56][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[56][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[56][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[56][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[56][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[56][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[56][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[56][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[56][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[56][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[56][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[56][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[56][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[56][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[56][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[56][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[56][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[56][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[56][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[56][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[56][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[56][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[56][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[56][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[56][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[56][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[56][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[56][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[56][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[56][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[56][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[56][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[56][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[56][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[56][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[56][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[56][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[56][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[56][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[56][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[56][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[56][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[56][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[56][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[56][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[56][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[56][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[56][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[56][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[56][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[56][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[56][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[56][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[56][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[56][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[56][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[56][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[56][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[56][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[56][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[56][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[56][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[56][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[56][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[56][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[56][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[56][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[56][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[56][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[56][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[56][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[56][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[56][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[56][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[56][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[56][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[56][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[56][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[56][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[56][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[56][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[56][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[56][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[56][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[56][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[56][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[56][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[56][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[56][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[56][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[56][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[56][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[56][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[56][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[56][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[56][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[56][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[56][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[56][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[56][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[56][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[56][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[56][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[56][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[56][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[56][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[56][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[56][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 56, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[56][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[56][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[56][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[56][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[56][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[56].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[56][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[57][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[57][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[57][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[57][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[57][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[57][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[57][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[57][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[57][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[57][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[57][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[57][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[57][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[57][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[57][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[57][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[57][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[57][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[57][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[57][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[57][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[57][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[57][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[57][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[57][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[57][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[57][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[57][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[57][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[57][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[57][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[57][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[57][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[57][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[57][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[57][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[57][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[57][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[57][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[57][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[57][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[57][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[57][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[57][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[57][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[57][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[57][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[57][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[57][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[57][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[57][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[57][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[57][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[57][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[57][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[57][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[57][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[57][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[57][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[57][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[57][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[57][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[57][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[57][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[57][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[57][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[57][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[57][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[57][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[57][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[57][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[57][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[57][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[57][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[57][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[57][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[57][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[57][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[57][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[57][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[57][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[57][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[57][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[57][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[57][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[57][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[57][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[57][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[57][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[57][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[57][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[57][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[57][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[57][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[57][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[57][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[57][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[57][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[57][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[57][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[57][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[57][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[57][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[57][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[57][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[57][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[57][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[57][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[57][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[57][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[57][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[57][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[57][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[57][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[57][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[57][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[57][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[57][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[57][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[57][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[57][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[57][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[57][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[57][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[57][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[57][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[57][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[57][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[57][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[57][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[57][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[57][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[57][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[57][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[57][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[57][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[57][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[57][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[57][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[57][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[57][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[57][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[57][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[57][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[57][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[57][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[57][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[57][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[57][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[57][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[57][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[57][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[57][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[57][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[57][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[57][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[57][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[57][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[57][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[57][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[57][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[57][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[57][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[57][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[57][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[57][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[57][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[57][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[57][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[57][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[57][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[57][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[57][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[57][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[57][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[57][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[57][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[57][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[57][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[57][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[57][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[57][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[57][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[57][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[57][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[57][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 57, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[57][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[57][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[57][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[57][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[57][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[57].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[57][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[58][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[58][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[58][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[58][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[58][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[58][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[58][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[58][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[58][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[58][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[58][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[58][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[58][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[58][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[58][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[58][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[58][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[58][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[58][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[58][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[58][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[58][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[58][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[58][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[58][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[58][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[58][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[58][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[58][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[58][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[58][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[58][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[58][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[58][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[58][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[58][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[58][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[58][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[58][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[58][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[58][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[58][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[58][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[58][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[58][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[58][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[58][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[58][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[58][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[58][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[58][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[58][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[58][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[58][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[58][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[58][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[58][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[58][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[58][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[58][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[58][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[58][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[58][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[58][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[58][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[58][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[58][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[58][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[58][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[58][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[58][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[58][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[58][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[58][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[58][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[58][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[58][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[58][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[58][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[58][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[58][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[58][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[58][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[58][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[58][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[58][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[58][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[58][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[58][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[58][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[58][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[58][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[58][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[58][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[58][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[58][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[58][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[58][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[58][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[58][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[58][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[58][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[58][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[58][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[58][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[58][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[58][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[58][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[58][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[58][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[58][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[58][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[58][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[58][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[58][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[58][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[58][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[58][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[58][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[58][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[58][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[58][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[58][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[58][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[58][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[58][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[58][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[58][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[58][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[58][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[58][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[58][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[58][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[58][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[58][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[58][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[58][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[58][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[58][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[58][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[58][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[58][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[58][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[58][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[58][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[58][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[58][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[58][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[58][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[58][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[58][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[58][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[58][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[58][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[58][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[58][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[58][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[58][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[58][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[58][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[58][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[58][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[58][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[58][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[58][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[58][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[58][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[58][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[58][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[58][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[58][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[58][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[58][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[58][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[58][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[58][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[58][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[58][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[58][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[58][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[58][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[58][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[58][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[58][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[58][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[58][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 58, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[58][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[58][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[58][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[58][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[58][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[58].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[58][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[59][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[59][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[59][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[59][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[59][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[59][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[59][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[59][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[59][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[59][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[59][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[59][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[59][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[59][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[59][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[59][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[59][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[59][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[59][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[59][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[59][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[59][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[59][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[59][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[59][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[59][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[59][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[59][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[59][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[59][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[59][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[59][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[59][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[59][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[59][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[59][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[59][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[59][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[59][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[59][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[59][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[59][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[59][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[59][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[59][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[59][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[59][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[59][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[59][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[59][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[59][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[59][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[59][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[59][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[59][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[59][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[59][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[59][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[59][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[59][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[59][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[59][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[59][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[59][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[59][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[59][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[59][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[59][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[59][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[59][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[59][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[59][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[59][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[59][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[59][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[59][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[59][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[59][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[59][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[59][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[59][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[59][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[59][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[59][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[59][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[59][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[59][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[59][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[59][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[59][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[59][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[59][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[59][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[59][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[59][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[59][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[59][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[59][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[59][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[59][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[59][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[59][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[59][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[59][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[59][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[59][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[59][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[59][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[59][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[59][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[59][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[59][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[59][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[59][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[59][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[59][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[59][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[59][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[59][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[59][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[59][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[59][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[59][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[59][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[59][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[59][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[59][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[59][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[59][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[59][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[59][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[59][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[59][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[59][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[59][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[59][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[59][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[59][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[59][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[59][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[59][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[59][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[59][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[59][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[59][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[59][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[59][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[59][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[59][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[59][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[59][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[59][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[59][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[59][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[59][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[59][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[59][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[59][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[59][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[59][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[59][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[59][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[59][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[59][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[59][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[59][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[59][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[59][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[59][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[59][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[59][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[59][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[59][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[59][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[59][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[59][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[59][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[59][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[59][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[59][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[59][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[59][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[59][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[59][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[59][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[59][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 59, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[59][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[59][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[59][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[59][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[59][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[59].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[59][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[60][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[60][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[60][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[60][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[60][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[60][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[60][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[60][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[60][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[60][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[60][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[60][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[60][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[60][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[60][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[60][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[60][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[60][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[60][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[60][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[60][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[60][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[60][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[60][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[60][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[60][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[60][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[60][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[60][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[60][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[60][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[60][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[60][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[60][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[60][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[60][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[60][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[60][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[60][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[60][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[60][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[60][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[60][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[60][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[60][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[60][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[60][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[60][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[60][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[60][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[60][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[60][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[60][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[60][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[60][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[60][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[60][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[60][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[60][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[60][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[60][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[60][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[60][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[60][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[60][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[60][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[60][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[60][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[60][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[60][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[60][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[60][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[60][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[60][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[60][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[60][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[60][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[60][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[60][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[60][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[60][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[60][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[60][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[60][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[60][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[60][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[60][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[60][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[60][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[60][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[60][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[60][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[60][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[60][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[60][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[60][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[60][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[60][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[60][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[60][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[60][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[60][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[60][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[60][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[60][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[60][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[60][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[60][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[60][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[60][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[60][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[60][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[60][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[60][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[60][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[60][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[60][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[60][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[60][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[60][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[60][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[60][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[60][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[60][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[60][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[60][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[60][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[60][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[60][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[60][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[60][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[60][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[60][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[60][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[60][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[60][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[60][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[60][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[60][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[60][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[60][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[60][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[60][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[60][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[60][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[60][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[60][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[60][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[60][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[60][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[60][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[60][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[60][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[60][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[60][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[60][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[60][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[60][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[60][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[60][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[60][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[60][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[60][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[60][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[60][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[60][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[60][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[60][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[60][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[60][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[60][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[60][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[60][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[60][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[60][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[60][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[60][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[60][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[60][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[60][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[60][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[60][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[60][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[60][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[60][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[60][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 60, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[60][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[60][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[60][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[60][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[60][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[60].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[60][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[61][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[61][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[61][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[61][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[61][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[61][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[61][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[61][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[61][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[61][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[61][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[61][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[61][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[61][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[61][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[61][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[61][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[61][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[61][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[61][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[61][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[61][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[61][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[61][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[61][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[61][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[61][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[61][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[61][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[61][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[61][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[61][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[61][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[61][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[61][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[61][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[61][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[61][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[61][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[61][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[61][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[61][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[61][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[61][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[61][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[61][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[61][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[61][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[61][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[61][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[61][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[61][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[61][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[61][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[61][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[61][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[61][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[61][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[61][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[61][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[61][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[61][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[61][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[61][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[61][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[61][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[61][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[61][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[61][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[61][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[61][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[61][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[61][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[61][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[61][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[61][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[61][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[61][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[61][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[61][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[61][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[61][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[61][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[61][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[61][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[61][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[61][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[61][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[61][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[61][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[61][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[61][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[61][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[61][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[61][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[61][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[61][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[61][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[61][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[61][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[61][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[61][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[61][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[61][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[61][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[61][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[61][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[61][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[61][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[61][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[61][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[61][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[61][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[61][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[61][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[61][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[61][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[61][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[61][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[61][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[61][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[61][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[61][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[61][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[61][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[61][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[61][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[61][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[61][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[61][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[61][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[61][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[61][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[61][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[61][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[61][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[61][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[61][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[61][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[61][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[61][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[61][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[61][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[61][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[61][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[61][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[61][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[61][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[61][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[61][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[61][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[61][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[61][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[61][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[61][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[61][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[61][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[61][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[61][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[61][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[61][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[61][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[61][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[61][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[61][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[61][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[61][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[61][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[61][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[61][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[61][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[61][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[61][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[61][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[61][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[61][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[61][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[61][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[61][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[61][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[61][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[61][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[61][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[61][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[61][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[61][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 61, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[61][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[61][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[61][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[61][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[61][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[61].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[61][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[62][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[62][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[62][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[62][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[62][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[62][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[62][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[62][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[62][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[62][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[62][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[62][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[62][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[62][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[62][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[62][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[62][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[62][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[62][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[62][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[62][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[62][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[62][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[62][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[62][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[62][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[62][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[62][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[62][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[62][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[62][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[62][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[62][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[62][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[62][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[62][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[62][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[62][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[62][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[62][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[62][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[62][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[62][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[62][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[62][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[62][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[62][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[62][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[62][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[62][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[62][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[62][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[62][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[62][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[62][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[62][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[62][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[62][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[62][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[62][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[62][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[62][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[62][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[62][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[62][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[62][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[62][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[62][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[62][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[62][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[62][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[62][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[62][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[62][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[62][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[62][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[62][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[62][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[62][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[62][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[62][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[62][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[62][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[62][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[62][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[62][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[62][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[62][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[62][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[62][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[62][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[62][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[62][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[62][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[62][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[62][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[62][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[62][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[62][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[62][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[62][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[62][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[62][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[62][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[62][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[62][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[62][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[62][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[62][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[62][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[62][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[62][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[62][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[62][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[62][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[62][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[62][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[62][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[62][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[62][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[62][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[62][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[62][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[62][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[62][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[62][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[62][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[62][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[62][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[62][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[62][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[62][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[62][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[62][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[62][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[62][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[62][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[62][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[62][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[62][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[62][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[62][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[62][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[62][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[62][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[62][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[62][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[62][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[62][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[62][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[62][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[62][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[62][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[62][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[62][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[62][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[62][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[62][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[62][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[62][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[62][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[62][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[62][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[62][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[62][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[62][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[62][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[62][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[62][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[62][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[62][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[62][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[62][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[62][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[62][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[62][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[62][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[62][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[62][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[62][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[62][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[62][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[62][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[62][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[62][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[62][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 62, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[62][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[62][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[62][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[62][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[62][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[62].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[62][31][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][0][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[63][0][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[63][0][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[63][0][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][0][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [0]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [0]  =   DownstreamStackBusLane[63][0][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [0]  =   DownstreamStackBusLane[63][0][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[0]  =   DownstreamStackBusLane[63][0][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][1][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[63][1][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[63][1][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[63][1][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][1][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [1]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [1]  =   DownstreamStackBusLane[63][1][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [1]  =   DownstreamStackBusLane[63][1][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[1]  =   DownstreamStackBusLane[63][1][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][2][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[63][2][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[63][2][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[63][2][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][2][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [2]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [2]  =   DownstreamStackBusLane[63][2][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [2]  =   DownstreamStackBusLane[63][2][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[2]  =   DownstreamStackBusLane[63][2][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][3][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[63][3][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[63][3][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[63][3][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][3][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [3]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [3]  =   DownstreamStackBusLane[63][3][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [3]  =   DownstreamStackBusLane[63][3][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[3]  =   DownstreamStackBusLane[63][3][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][4][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[63][4][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[63][4][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[63][4][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][4][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [4]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [4]  =   DownstreamStackBusLane[63][4][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [4]  =   DownstreamStackBusLane[63][4][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[4]  =   DownstreamStackBusLane[63][4][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][5][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[63][5][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[63][5][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[63][5][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][5][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [5]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [5]  =   DownstreamStackBusLane[63][5][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [5]  =   DownstreamStackBusLane[63][5][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[5]  =   DownstreamStackBusLane[63][5][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][6][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[63][6][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[63][6][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[63][6][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][6][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [6]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [6]  =   DownstreamStackBusLane[63][6][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [6]  =   DownstreamStackBusLane[63][6][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[6]  =   DownstreamStackBusLane[63][6][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][7][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[63][7][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[63][7][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[63][7][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][7][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [7]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [7]  =   DownstreamStackBusLane[63][7][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [7]  =   DownstreamStackBusLane[63][7][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[7]  =   DownstreamStackBusLane[63][7][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][8][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[63][8][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[63][8][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[63][8][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][8][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [8]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [8]  =   DownstreamStackBusLane[63][8][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [8]  =   DownstreamStackBusLane[63][8][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[8]  =   DownstreamStackBusLane[63][8][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][9][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[63][9][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[63][9][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[63][9][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][9][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [9]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [9]  =   DownstreamStackBusLane[63][9][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [9]  =   DownstreamStackBusLane[63][9][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[9]  =   DownstreamStackBusLane[63][9][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][10][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[63][10][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[63][10][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[63][10][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][10][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [10]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [10]  =   DownstreamStackBusLane[63][10][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [10]  =   DownstreamStackBusLane[63][10][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[10]  =   DownstreamStackBusLane[63][10][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][11][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[63][11][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[63][11][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[63][11][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][11][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [11]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [11]  =   DownstreamStackBusLane[63][11][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [11]  =   DownstreamStackBusLane[63][11][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[11]  =   DownstreamStackBusLane[63][11][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][12][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[63][12][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[63][12][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[63][12][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][12][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [12]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [12]  =   DownstreamStackBusLane[63][12][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [12]  =   DownstreamStackBusLane[63][12][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[12]  =   DownstreamStackBusLane[63][12][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][13][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[63][13][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[63][13][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[63][13][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][13][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [13]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [13]  =   DownstreamStackBusLane[63][13][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [13]  =   DownstreamStackBusLane[63][13][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[13]  =   DownstreamStackBusLane[63][13][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][14][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[63][14][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[63][14][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[63][14][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][14][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [14]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [14]  =   DownstreamStackBusLane[63][14][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [14]  =   DownstreamStackBusLane[63][14][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[14]  =   DownstreamStackBusLane[63][14][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][15][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[63][15][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[63][15][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[63][15][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][15][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [15]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [15]  =   DownstreamStackBusLane[63][15][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [15]  =   DownstreamStackBusLane[63][15][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[15]  =   DownstreamStackBusLane[63][15][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][16][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[63][16][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[63][16][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[63][16][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][16][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [16]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [16]  =   DownstreamStackBusLane[63][16][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [16]  =   DownstreamStackBusLane[63][16][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[16]  =   DownstreamStackBusLane[63][16][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][17][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[63][17][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[63][17][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[63][17][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][17][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [17]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [17]  =   DownstreamStackBusLane[63][17][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [17]  =   DownstreamStackBusLane[63][17][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[17]  =   DownstreamStackBusLane[63][17][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][18][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[63][18][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[63][18][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[63][18][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][18][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [18]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [18]  =   DownstreamStackBusLane[63][18][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [18]  =   DownstreamStackBusLane[63][18][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[18]  =   DownstreamStackBusLane[63][18][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][19][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[63][19][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[63][19][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[63][19][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][19][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [19]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [19]  =   DownstreamStackBusLane[63][19][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [19]  =   DownstreamStackBusLane[63][19][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[19]  =   DownstreamStackBusLane[63][19][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][20][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[63][20][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[63][20][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[63][20][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][20][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [20]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [20]  =   DownstreamStackBusLane[63][20][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [20]  =   DownstreamStackBusLane[63][20][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[20]  =   DownstreamStackBusLane[63][20][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][21][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[63][21][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[63][21][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[63][21][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][21][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [21]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [21]  =   DownstreamStackBusLane[63][21][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [21]  =   DownstreamStackBusLane[63][21][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[21]  =   DownstreamStackBusLane[63][21][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][22][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[63][22][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[63][22][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[63][22][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][22][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [22]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [22]  =   DownstreamStackBusLane[63][22][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [22]  =   DownstreamStackBusLane[63][22][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[22]  =   DownstreamStackBusLane[63][22][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][23][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[63][23][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[63][23][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[63][23][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][23][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [23]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [23]  =   DownstreamStackBusLane[63][23][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [23]  =   DownstreamStackBusLane[63][23][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[23]  =   DownstreamStackBusLane[63][23][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][24][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[63][24][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[63][24][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[63][24][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][24][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [24]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [24]  =   DownstreamStackBusLane[63][24][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [24]  =   DownstreamStackBusLane[63][24][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[24]  =   DownstreamStackBusLane[63][24][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][25][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[63][25][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[63][25][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[63][25][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][25][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [25]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [25]  =   DownstreamStackBusLane[63][25][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [25]  =   DownstreamStackBusLane[63][25][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[25]  =   DownstreamStackBusLane[63][25][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][26][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[63][26][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[63][26][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[63][26][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][26][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [26]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [26]  =   DownstreamStackBusLane[63][26][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [26]  =   DownstreamStackBusLane[63][26][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[26]  =   DownstreamStackBusLane[63][26][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][27][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[63][27][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[63][27][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[63][27][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][27][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [27]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [27]  =   DownstreamStackBusLane[63][27][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [27]  =   DownstreamStackBusLane[63][27][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[27]  =   DownstreamStackBusLane[63][27][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][28][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[63][28][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[63][28][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[63][28][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][28][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [28]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [28]  =   DownstreamStackBusLane[63][28][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [28]  =   DownstreamStackBusLane[63][28][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[28]  =   DownstreamStackBusLane[63][28][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][29][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[63][29][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[63][29][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[63][29][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][29][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [29]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [29]  =   DownstreamStackBusLane[63][29][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [29]  =   DownstreamStackBusLane[63][29][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[29]  =   DownstreamStackBusLane[63][29][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][30][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[63][30][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[63][30][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[63][30][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][30][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [30]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [30]  =   DownstreamStackBusLane[63][30][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [30]  =   DownstreamStackBusLane[63][30][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[30]  =   DownstreamStackBusLane[63][30][1].std__pe__lane_strm_data_valid ;
          end
        
        // PE 63, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][31][0].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[63][31][0].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[63][31][0].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[0].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[63][31][0].std__pe__lane_strm_data_valid ;
          end
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][31][1].pe__std__lane_strm_ready   =   system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.std__mrc__lane_ready [31]    ;
        always @(*)
          begin
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_cntl_e1 [31]  =   DownstreamStackBusLane[63][31][1].std__pe__lane_strm_cntl       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_data_e1 [31]  =   DownstreamStackBusLane[63][31][1].std__pe__lane_strm_data       ;
            system_inst.manager_array_inst.mgr_inst[63].manager.mrc_cntl_strm_inst[1].mrc_cntl.mrc__std__lane_valid_e1[31]  =   DownstreamStackBusLane[63][31][1].std__pe__lane_strm_data_valid ;
          end
        