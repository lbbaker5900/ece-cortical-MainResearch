
  // General control and status                                                
  wire                                        sys__pe0__allSynchronized     ;
  wire                                        pe0__sys__thisSynchronized    ;
  wire                                        pe0__sys__ready               ;
  wire                                        pe0__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe1__allSynchronized     ;
  wire                                        pe1__sys__thisSynchronized    ;
  wire                                        pe1__sys__ready               ;
  wire                                        pe1__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe2__allSynchronized     ;
  wire                                        pe2__sys__thisSynchronized    ;
  wire                                        pe2__sys__ready               ;
  wire                                        pe2__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe3__allSynchronized     ;
  wire                                        pe3__sys__thisSynchronized    ;
  wire                                        pe3__sys__ready               ;
  wire                                        pe3__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe4__allSynchronized     ;
  wire                                        pe4__sys__thisSynchronized    ;
  wire                                        pe4__sys__ready               ;
  wire                                        pe4__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe5__allSynchronized     ;
  wire                                        pe5__sys__thisSynchronized    ;
  wire                                        pe5__sys__ready               ;
  wire                                        pe5__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe6__allSynchronized     ;
  wire                                        pe6__sys__thisSynchronized    ;
  wire                                        pe6__sys__ready               ;
  wire                                        pe6__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe7__allSynchronized     ;
  wire                                        pe7__sys__thisSynchronized    ;
  wire                                        pe7__sys__ready               ;
  wire                                        pe7__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe8__allSynchronized     ;
  wire                                        pe8__sys__thisSynchronized    ;
  wire                                        pe8__sys__ready               ;
  wire                                        pe8__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe9__allSynchronized     ;
  wire                                        pe9__sys__thisSynchronized    ;
  wire                                        pe9__sys__ready               ;
  wire                                        pe9__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe10__allSynchronized     ;
  wire                                        pe10__sys__thisSynchronized    ;
  wire                                        pe10__sys__ready               ;
  wire                                        pe10__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe11__allSynchronized     ;
  wire                                        pe11__sys__thisSynchronized    ;
  wire                                        pe11__sys__ready               ;
  wire                                        pe11__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe12__allSynchronized     ;
  wire                                        pe12__sys__thisSynchronized    ;
  wire                                        pe12__sys__ready               ;
  wire                                        pe12__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe13__allSynchronized     ;
  wire                                        pe13__sys__thisSynchronized    ;
  wire                                        pe13__sys__ready               ;
  wire                                        pe13__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe14__allSynchronized     ;
  wire                                        pe14__sys__thisSynchronized    ;
  wire                                        pe14__sys__ready               ;
  wire                                        pe14__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe15__allSynchronized     ;
  wire                                        pe15__sys__thisSynchronized    ;
  wire                                        pe15__sys__ready               ;
  wire                                        pe15__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe16__allSynchronized     ;
  wire                                        pe16__sys__thisSynchronized    ;
  wire                                        pe16__sys__ready               ;
  wire                                        pe16__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe17__allSynchronized     ;
  wire                                        pe17__sys__thisSynchronized    ;
  wire                                        pe17__sys__ready               ;
  wire                                        pe17__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe18__allSynchronized     ;
  wire                                        pe18__sys__thisSynchronized    ;
  wire                                        pe18__sys__ready               ;
  wire                                        pe18__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe19__allSynchronized     ;
  wire                                        pe19__sys__thisSynchronized    ;
  wire                                        pe19__sys__ready               ;
  wire                                        pe19__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe20__allSynchronized     ;
  wire                                        pe20__sys__thisSynchronized    ;
  wire                                        pe20__sys__ready               ;
  wire                                        pe20__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe21__allSynchronized     ;
  wire                                        pe21__sys__thisSynchronized    ;
  wire                                        pe21__sys__ready               ;
  wire                                        pe21__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe22__allSynchronized     ;
  wire                                        pe22__sys__thisSynchronized    ;
  wire                                        pe22__sys__ready               ;
  wire                                        pe22__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe23__allSynchronized     ;
  wire                                        pe23__sys__thisSynchronized    ;
  wire                                        pe23__sys__ready               ;
  wire                                        pe23__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe24__allSynchronized     ;
  wire                                        pe24__sys__thisSynchronized    ;
  wire                                        pe24__sys__ready               ;
  wire                                        pe24__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe25__allSynchronized     ;
  wire                                        pe25__sys__thisSynchronized    ;
  wire                                        pe25__sys__ready               ;
  wire                                        pe25__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe26__allSynchronized     ;
  wire                                        pe26__sys__thisSynchronized    ;
  wire                                        pe26__sys__ready               ;
  wire                                        pe26__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe27__allSynchronized     ;
  wire                                        pe27__sys__thisSynchronized    ;
  wire                                        pe27__sys__ready               ;
  wire                                        pe27__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe28__allSynchronized     ;
  wire                                        pe28__sys__thisSynchronized    ;
  wire                                        pe28__sys__ready               ;
  wire                                        pe28__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe29__allSynchronized     ;
  wire                                        pe29__sys__thisSynchronized    ;
  wire                                        pe29__sys__ready               ;
  wire                                        pe29__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe30__allSynchronized     ;
  wire                                        pe30__sys__thisSynchronized    ;
  wire                                        pe30__sys__ready               ;
  wire                                        pe30__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe31__allSynchronized     ;
  wire                                        pe31__sys__thisSynchronized    ;
  wire                                        pe31__sys__ready               ;
  wire                                        pe31__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe32__allSynchronized     ;
  wire                                        pe32__sys__thisSynchronized    ;
  wire                                        pe32__sys__ready               ;
  wire                                        pe32__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe33__allSynchronized     ;
  wire                                        pe33__sys__thisSynchronized    ;
  wire                                        pe33__sys__ready               ;
  wire                                        pe33__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe34__allSynchronized     ;
  wire                                        pe34__sys__thisSynchronized    ;
  wire                                        pe34__sys__ready               ;
  wire                                        pe34__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe35__allSynchronized     ;
  wire                                        pe35__sys__thisSynchronized    ;
  wire                                        pe35__sys__ready               ;
  wire                                        pe35__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe36__allSynchronized     ;
  wire                                        pe36__sys__thisSynchronized    ;
  wire                                        pe36__sys__ready               ;
  wire                                        pe36__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe37__allSynchronized     ;
  wire                                        pe37__sys__thisSynchronized    ;
  wire                                        pe37__sys__ready               ;
  wire                                        pe37__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe38__allSynchronized     ;
  wire                                        pe38__sys__thisSynchronized    ;
  wire                                        pe38__sys__ready               ;
  wire                                        pe38__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe39__allSynchronized     ;
  wire                                        pe39__sys__thisSynchronized    ;
  wire                                        pe39__sys__ready               ;
  wire                                        pe39__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe40__allSynchronized     ;
  wire                                        pe40__sys__thisSynchronized    ;
  wire                                        pe40__sys__ready               ;
  wire                                        pe40__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe41__allSynchronized     ;
  wire                                        pe41__sys__thisSynchronized    ;
  wire                                        pe41__sys__ready               ;
  wire                                        pe41__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe42__allSynchronized     ;
  wire                                        pe42__sys__thisSynchronized    ;
  wire                                        pe42__sys__ready               ;
  wire                                        pe42__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe43__allSynchronized     ;
  wire                                        pe43__sys__thisSynchronized    ;
  wire                                        pe43__sys__ready               ;
  wire                                        pe43__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe44__allSynchronized     ;
  wire                                        pe44__sys__thisSynchronized    ;
  wire                                        pe44__sys__ready               ;
  wire                                        pe44__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe45__allSynchronized     ;
  wire                                        pe45__sys__thisSynchronized    ;
  wire                                        pe45__sys__ready               ;
  wire                                        pe45__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe46__allSynchronized     ;
  wire                                        pe46__sys__thisSynchronized    ;
  wire                                        pe46__sys__ready               ;
  wire                                        pe46__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe47__allSynchronized     ;
  wire                                        pe47__sys__thisSynchronized    ;
  wire                                        pe47__sys__ready               ;
  wire                                        pe47__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe48__allSynchronized     ;
  wire                                        pe48__sys__thisSynchronized    ;
  wire                                        pe48__sys__ready               ;
  wire                                        pe48__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe49__allSynchronized     ;
  wire                                        pe49__sys__thisSynchronized    ;
  wire                                        pe49__sys__ready               ;
  wire                                        pe49__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe50__allSynchronized     ;
  wire                                        pe50__sys__thisSynchronized    ;
  wire                                        pe50__sys__ready               ;
  wire                                        pe50__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe51__allSynchronized     ;
  wire                                        pe51__sys__thisSynchronized    ;
  wire                                        pe51__sys__ready               ;
  wire                                        pe51__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe52__allSynchronized     ;
  wire                                        pe52__sys__thisSynchronized    ;
  wire                                        pe52__sys__ready               ;
  wire                                        pe52__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe53__allSynchronized     ;
  wire                                        pe53__sys__thisSynchronized    ;
  wire                                        pe53__sys__ready               ;
  wire                                        pe53__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe54__allSynchronized     ;
  wire                                        pe54__sys__thisSynchronized    ;
  wire                                        pe54__sys__ready               ;
  wire                                        pe54__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe55__allSynchronized     ;
  wire                                        pe55__sys__thisSynchronized    ;
  wire                                        pe55__sys__ready               ;
  wire                                        pe55__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe56__allSynchronized     ;
  wire                                        pe56__sys__thisSynchronized    ;
  wire                                        pe56__sys__ready               ;
  wire                                        pe56__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe57__allSynchronized     ;
  wire                                        pe57__sys__thisSynchronized    ;
  wire                                        pe57__sys__ready               ;
  wire                                        pe57__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe58__allSynchronized     ;
  wire                                        pe58__sys__thisSynchronized    ;
  wire                                        pe58__sys__ready               ;
  wire                                        pe58__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe59__allSynchronized     ;
  wire                                        pe59__sys__thisSynchronized    ;
  wire                                        pe59__sys__ready               ;
  wire                                        pe59__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe60__allSynchronized     ;
  wire                                        pe60__sys__thisSynchronized    ;
  wire                                        pe60__sys__ready               ;
  wire                                        pe60__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe61__allSynchronized     ;
  wire                                        pe61__sys__thisSynchronized    ;
  wire                                        pe61__sys__ready               ;
  wire                                        pe61__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe62__allSynchronized     ;
  wire                                        pe62__sys__thisSynchronized    ;
  wire                                        pe62__sys__ready               ;
  wire                                        pe62__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe63__allSynchronized     ;
  wire                                        pe63__sys__thisSynchronized    ;
  wire                                        pe63__sys__ready               ;
  wire                                        pe63__sys__complete            ;