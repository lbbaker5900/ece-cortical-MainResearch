

  // Convert the mgrId of the pointer to a bit mask
  always @(*)
    begin
      case(currPtrManager)
      6'd0 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000000000000000000001  ; 
        end
      6'd1 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000000000000000000010  ; 
        end
      6'd2 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000000000000000000100  ; 
        end
      6'd3 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000000000000000001000  ; 
        end
      6'd4 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000000000000000010000  ; 
        end
      6'd5 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000000000000000100000  ; 
        end
      6'd6 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000000000000001000000  ; 
        end
      6'd7 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000000000000010000000  ; 
        end
      6'd8 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000000000000100000000  ; 
        end
      6'd9 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000000000001000000000  ; 
        end
      6'd10 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000000000010000000000  ; 
        end
      6'd11 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000000000100000000000  ; 
        end
      6'd12 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000000001000000000000  ; 
        end
      6'd13 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000000010000000000000  ; 
        end
      6'd14 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000000100000000000000  ; 
        end
      6'd15 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000001000000000000000  ; 
        end
      6'd16 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000010000000000000000  ; 
        end
      6'd17 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000000100000000000000000  ; 
        end
      6'd18 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000001000000000000000000  ; 
        end
      6'd19 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000010000000000000000000  ; 
        end
      6'd20 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000000100000000000000000000  ; 
        end
      6'd21 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000001000000000000000000000  ; 
        end
      6'd22 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000010000000000000000000000  ; 
        end
      6'd23 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000000100000000000000000000000  ; 
        end
      6'd24 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000001000000000000000000000000  ; 
        end
      6'd25 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000010000000000000000000000000  ; 
        end
      6'd26 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000000100000000000000000000000000  ; 
        end
      6'd27 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000001000000000000000000000000000  ; 
        end
      6'd28 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000010000000000000000000000000000  ; 
        end
      6'd29 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000000100000000000000000000000000000  ; 
        end
      6'd30 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000001000000000000000000000000000000  ; 
        end
      6'd31 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000010000000000000000000000000000000  ; 
        end
      6'd32 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000000100000000000000000000000000000000  ; 
        end
      6'd33 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000001000000000000000000000000000000000  ; 
        end
      6'd34 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000010000000000000000000000000000000000  ; 
        end
      6'd35 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000000100000000000000000000000000000000000  ; 
        end
      6'd36 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000001000000000000000000000000000000000000  ; 
        end
      6'd37 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000010000000000000000000000000000000000000  ; 
        end
      6'd38 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000000100000000000000000000000000000000000000  ; 
        end
      6'd39 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000001000000000000000000000000000000000000000  ; 
        end
      6'd40 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000010000000000000000000000000000000000000000  ; 
        end
      6'd41 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000000100000000000000000000000000000000000000000  ; 
        end
      6'd42 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000001000000000000000000000000000000000000000000  ; 
        end
      6'd43 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000010000000000000000000000000000000000000000000  ; 
        end
      6'd44 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000000100000000000000000000000000000000000000000000  ; 
        end
      6'd45 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000001000000000000000000000000000000000000000000000  ; 
        end
      6'd46 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000010000000000000000000000000000000000000000000000  ; 
        end
      6'd47 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000000100000000000000000000000000000000000000000000000  ; 
        end
      6'd48 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000001000000000000000000000000000000000000000000000000  ; 
        end
      6'd49 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000010000000000000000000000000000000000000000000000000  ; 
        end
      6'd50 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000000100000000000000000000000000000000000000000000000000  ; 
        end
      6'd51 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000001000000000000000000000000000000000000000000000000000  ; 
        end
      6'd52 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000010000000000000000000000000000000000000000000000000000  ; 
        end
      6'd53 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000000100000000000000000000000000000000000000000000000000000  ; 
        end
      6'd54 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000001000000000000000000000000000000000000000000000000000000  ; 
        end
      6'd55 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000010000000000000000000000000000000000000000000000000000000  ; 
        end
      6'd56 :
        begin
          currPtrDestBitMaskAddr = 64'b0000000100000000000000000000000000000000000000000000000000000000  ; 
        end
      6'd57 :
        begin
          currPtrDestBitMaskAddr = 64'b0000001000000000000000000000000000000000000000000000000000000000  ; 
        end
      6'd58 :
        begin
          currPtrDestBitMaskAddr = 64'b0000010000000000000000000000000000000000000000000000000000000000  ; 
        end
      6'd59 :
        begin
          currPtrDestBitMaskAddr = 64'b0000100000000000000000000000000000000000000000000000000000000000  ; 
        end
      6'd60 :
        begin
          currPtrDestBitMaskAddr = 64'b0001000000000000000000000000000000000000000000000000000000000000  ; 
        end
      6'd61 :
        begin
          currPtrDestBitMaskAddr = 64'b0010000000000000000000000000000000000000000000000000000000000000  ; 
        end
      6'd62 :
        begin
          currPtrDestBitMaskAddr = 64'b0100000000000000000000000000000000000000000000000000000000000000  ; 
        end
      6'd63 :
        begin
          currPtrDestBitMaskAddr = 64'b1000000000000000000000000000000000000000000000000000000000000000  ; 
        end
      default:
        begin
          currPtrDestBitMaskAddr = 64'd0 ; 
        end
      endcase
    end
