`ifndef _sd_memory_vh
`define _sd_memory_vh

/*****************************************************************

    File name   : sd_memory.vh
    Author      : Lee Baker
    Affiliation : North Carolina State University, Raleigh, NC
    Date        : Mar 2017
    email       : lbbaker@ncsu.edu

*****************************************************************/


//--------------------------------------------------------
  
//------------------------------------------------------------------------------------------------------------


`endif
