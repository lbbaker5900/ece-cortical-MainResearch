
   reg [`MGR_MGR_ID_BITMASK_RANGE      ] thisMgrBitMask       ; 