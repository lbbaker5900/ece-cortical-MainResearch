
  // General control and status                                                
  wire                                        sys__pe0__allSynchronized     ;
  wire                                        pe0__sys__thisSynchronized    ;
  wire                                        pe0__sys__ready               ;
  wire                                        pe0__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe1__allSynchronized     ;
  wire                                        pe1__sys__thisSynchronized    ;
  wire                                        pe1__sys__ready               ;
  wire                                        pe1__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe2__allSynchronized     ;
  wire                                        pe2__sys__thisSynchronized    ;
  wire                                        pe2__sys__ready               ;
  wire                                        pe2__sys__complete            ;
  // General control and status                                                
  wire                                        sys__pe3__allSynchronized     ;
  wire                                        pe3__sys__thisSynchronized    ;
  wire                                        pe3__sys__ready               ;
  wire                                        pe3__sys__complete            ;