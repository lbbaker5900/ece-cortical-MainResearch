
 assign    stu__mgr0__valid       =    pe0__stu__valid          ;
 assign    stu__mgr0__cntl        =    pe0__stu__cntl           ;
 assign    stu__pe0__ready        =    mgr0__stu__ready         ;
 assign    stu__mgr0__type        =    pe0__stu__type           ;
 assign    stu__mgr0__data        =    pe0__stu__data           ;
 assign    stu__mgr0__oob_data    =    pe0__stu__oob_data       ;

 assign    stu__mgr1__valid       =    pe1__stu__valid          ;
 assign    stu__mgr1__cntl        =    pe1__stu__cntl           ;
 assign    stu__pe1__ready        =    mgr1__stu__ready         ;
 assign    stu__mgr1__type        =    pe1__stu__type           ;
 assign    stu__mgr1__data        =    pe1__stu__data           ;
 assign    stu__mgr1__oob_data    =    pe1__stu__oob_data       ;

 assign    stu__mgr2__valid       =    pe2__stu__valid          ;
 assign    stu__mgr2__cntl        =    pe2__stu__cntl           ;
 assign    stu__pe2__ready        =    mgr2__stu__ready         ;
 assign    stu__mgr2__type        =    pe2__stu__type           ;
 assign    stu__mgr2__data        =    pe2__stu__data           ;
 assign    stu__mgr2__oob_data    =    pe2__stu__oob_data       ;

 assign    stu__mgr3__valid       =    pe3__stu__valid          ;
 assign    stu__mgr3__cntl        =    pe3__stu__cntl           ;
 assign    stu__pe3__ready        =    mgr3__stu__ready         ;
 assign    stu__mgr3__type        =    pe3__stu__type           ;
 assign    stu__mgr3__data        =    pe3__stu__data           ;
 assign    stu__mgr3__oob_data    =    pe3__stu__oob_data       ;

