
        begin
          forever
            begin
              // Observe NoC packets sent from manager 0
              @(vLocalToNoC[0].cb_p);
              if ((vLocalToNoC[0].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[0].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 0);
                  local_noc_pkt_sent [0] = new();
                  local_noc_pkt_sent [0].header_destination_address  = vLocalToNoC[0].locl__noc__dp_data     ;
                  local_noc_pkt_sent [0].header_source               = 0                                     ;
                  local_noc_pkt_sent [0].header_address_type         = vLocalToNoC[0].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [0].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [0].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 0, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [0]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 1
              @(vLocalToNoC[1].cb_p);
              if ((vLocalToNoC[1].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[1].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 1);
                  local_noc_pkt_sent [1] = new();
                  local_noc_pkt_sent [1].header_destination_address  = vLocalToNoC[1].locl__noc__dp_data     ;
                  local_noc_pkt_sent [1].header_source               = 1                                     ;
                  local_noc_pkt_sent [1].header_address_type         = vLocalToNoC[1].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [1].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [1].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 1, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [1]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 2
              @(vLocalToNoC[2].cb_p);
              if ((vLocalToNoC[2].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[2].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 2);
                  local_noc_pkt_sent [2] = new();
                  local_noc_pkt_sent [2].header_destination_address  = vLocalToNoC[2].locl__noc__dp_data     ;
                  local_noc_pkt_sent [2].header_source               = 2                                     ;
                  local_noc_pkt_sent [2].header_address_type         = vLocalToNoC[2].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [2].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [2].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 2, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [2]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 3
              @(vLocalToNoC[3].cb_p);
              if ((vLocalToNoC[3].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[3].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 3);
                  local_noc_pkt_sent [3] = new();
                  local_noc_pkt_sent [3].header_destination_address  = vLocalToNoC[3].locl__noc__dp_data     ;
                  local_noc_pkt_sent [3].header_source               = 3                                     ;
                  local_noc_pkt_sent [3].header_address_type         = vLocalToNoC[3].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [3].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [3].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 3, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [3]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 4
              @(vLocalToNoC[4].cb_p);
              if ((vLocalToNoC[4].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[4].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 4);
                  local_noc_pkt_sent [4] = new();
                  local_noc_pkt_sent [4].header_destination_address  = vLocalToNoC[4].locl__noc__dp_data     ;
                  local_noc_pkt_sent [4].header_source               = 4                                     ;
                  local_noc_pkt_sent [4].header_address_type         = vLocalToNoC[4].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [4].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [4].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 4, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [4]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 5
              @(vLocalToNoC[5].cb_p);
              if ((vLocalToNoC[5].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[5].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 5);
                  local_noc_pkt_sent [5] = new();
                  local_noc_pkt_sent [5].header_destination_address  = vLocalToNoC[5].locl__noc__dp_data     ;
                  local_noc_pkt_sent [5].header_source               = 5                                     ;
                  local_noc_pkt_sent [5].header_address_type         = vLocalToNoC[5].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [5].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [5].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 5, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [5]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 6
              @(vLocalToNoC[6].cb_p);
              if ((vLocalToNoC[6].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[6].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 6);
                  local_noc_pkt_sent [6] = new();
                  local_noc_pkt_sent [6].header_destination_address  = vLocalToNoC[6].locl__noc__dp_data     ;
                  local_noc_pkt_sent [6].header_source               = 6                                     ;
                  local_noc_pkt_sent [6].header_address_type         = vLocalToNoC[6].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [6].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [6].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 6, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [6]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 7
              @(vLocalToNoC[7].cb_p);
              if ((vLocalToNoC[7].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[7].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 7);
                  local_noc_pkt_sent [7] = new();
                  local_noc_pkt_sent [7].header_destination_address  = vLocalToNoC[7].locl__noc__dp_data     ;
                  local_noc_pkt_sent [7].header_source               = 7                                     ;
                  local_noc_pkt_sent [7].header_address_type         = vLocalToNoC[7].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [7].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [7].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 7, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [7]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 8
              @(vLocalToNoC[8].cb_p);
              if ((vLocalToNoC[8].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[8].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 8);
                  local_noc_pkt_sent [8] = new();
                  local_noc_pkt_sent [8].header_destination_address  = vLocalToNoC[8].locl__noc__dp_data     ;
                  local_noc_pkt_sent [8].header_source               = 8                                     ;
                  local_noc_pkt_sent [8].header_address_type         = vLocalToNoC[8].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [8].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [8].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 8, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [8]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 9
              @(vLocalToNoC[9].cb_p);
              if ((vLocalToNoC[9].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[9].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 9);
                  local_noc_pkt_sent [9] = new();
                  local_noc_pkt_sent [9].header_destination_address  = vLocalToNoC[9].locl__noc__dp_data     ;
                  local_noc_pkt_sent [9].header_source               = 9                                     ;
                  local_noc_pkt_sent [9].header_address_type         = vLocalToNoC[9].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [9].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [9].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 9, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [9]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 10
              @(vLocalToNoC[10].cb_p);
              if ((vLocalToNoC[10].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[10].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 10);
                  local_noc_pkt_sent [10] = new();
                  local_noc_pkt_sent [10].header_destination_address  = vLocalToNoC[10].locl__noc__dp_data     ;
                  local_noc_pkt_sent [10].header_source               = 10                                     ;
                  local_noc_pkt_sent [10].header_address_type         = vLocalToNoC[10].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [10].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [10].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 10, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [10]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 11
              @(vLocalToNoC[11].cb_p);
              if ((vLocalToNoC[11].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[11].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 11);
                  local_noc_pkt_sent [11] = new();
                  local_noc_pkt_sent [11].header_destination_address  = vLocalToNoC[11].locl__noc__dp_data     ;
                  local_noc_pkt_sent [11].header_source               = 11                                     ;
                  local_noc_pkt_sent [11].header_address_type         = vLocalToNoC[11].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [11].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [11].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 11, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [11]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 12
              @(vLocalToNoC[12].cb_p);
              if ((vLocalToNoC[12].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[12].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 12);
                  local_noc_pkt_sent [12] = new();
                  local_noc_pkt_sent [12].header_destination_address  = vLocalToNoC[12].locl__noc__dp_data     ;
                  local_noc_pkt_sent [12].header_source               = 12                                     ;
                  local_noc_pkt_sent [12].header_address_type         = vLocalToNoC[12].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [12].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [12].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 12, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [12]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 13
              @(vLocalToNoC[13].cb_p);
              if ((vLocalToNoC[13].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[13].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 13);
                  local_noc_pkt_sent [13] = new();
                  local_noc_pkt_sent [13].header_destination_address  = vLocalToNoC[13].locl__noc__dp_data     ;
                  local_noc_pkt_sent [13].header_source               = 13                                     ;
                  local_noc_pkt_sent [13].header_address_type         = vLocalToNoC[13].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [13].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [13].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 13, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [13]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 14
              @(vLocalToNoC[14].cb_p);
              if ((vLocalToNoC[14].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[14].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 14);
                  local_noc_pkt_sent [14] = new();
                  local_noc_pkt_sent [14].header_destination_address  = vLocalToNoC[14].locl__noc__dp_data     ;
                  local_noc_pkt_sent [14].header_source               = 14                                     ;
                  local_noc_pkt_sent [14].header_address_type         = vLocalToNoC[14].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [14].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [14].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 14, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [14]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 15
              @(vLocalToNoC[15].cb_p);
              if ((vLocalToNoC[15].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[15].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 15);
                  local_noc_pkt_sent [15] = new();
                  local_noc_pkt_sent [15].header_destination_address  = vLocalToNoC[15].locl__noc__dp_data     ;
                  local_noc_pkt_sent [15].header_source               = 15                                     ;
                  local_noc_pkt_sent [15].header_address_type         = vLocalToNoC[15].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [15].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [15].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 15, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [15]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 16
              @(vLocalToNoC[16].cb_p);
              if ((vLocalToNoC[16].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[16].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 16);
                  local_noc_pkt_sent [16] = new();
                  local_noc_pkt_sent [16].header_destination_address  = vLocalToNoC[16].locl__noc__dp_data     ;
                  local_noc_pkt_sent [16].header_source               = 16                                     ;
                  local_noc_pkt_sent [16].header_address_type         = vLocalToNoC[16].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [16].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [16].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 16, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [16]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 17
              @(vLocalToNoC[17].cb_p);
              if ((vLocalToNoC[17].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[17].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 17);
                  local_noc_pkt_sent [17] = new();
                  local_noc_pkt_sent [17].header_destination_address  = vLocalToNoC[17].locl__noc__dp_data     ;
                  local_noc_pkt_sent [17].header_source               = 17                                     ;
                  local_noc_pkt_sent [17].header_address_type         = vLocalToNoC[17].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [17].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [17].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 17, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [17]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 18
              @(vLocalToNoC[18].cb_p);
              if ((vLocalToNoC[18].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[18].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 18);
                  local_noc_pkt_sent [18] = new();
                  local_noc_pkt_sent [18].header_destination_address  = vLocalToNoC[18].locl__noc__dp_data     ;
                  local_noc_pkt_sent [18].header_source               = 18                                     ;
                  local_noc_pkt_sent [18].header_address_type         = vLocalToNoC[18].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [18].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [18].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 18, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [18]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 19
              @(vLocalToNoC[19].cb_p);
              if ((vLocalToNoC[19].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[19].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 19);
                  local_noc_pkt_sent [19] = new();
                  local_noc_pkt_sent [19].header_destination_address  = vLocalToNoC[19].locl__noc__dp_data     ;
                  local_noc_pkt_sent [19].header_source               = 19                                     ;
                  local_noc_pkt_sent [19].header_address_type         = vLocalToNoC[19].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [19].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [19].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 19, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [19]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 20
              @(vLocalToNoC[20].cb_p);
              if ((vLocalToNoC[20].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[20].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 20);
                  local_noc_pkt_sent [20] = new();
                  local_noc_pkt_sent [20].header_destination_address  = vLocalToNoC[20].locl__noc__dp_data     ;
                  local_noc_pkt_sent [20].header_source               = 20                                     ;
                  local_noc_pkt_sent [20].header_address_type         = vLocalToNoC[20].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [20].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [20].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 20, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [20]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 21
              @(vLocalToNoC[21].cb_p);
              if ((vLocalToNoC[21].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[21].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 21);
                  local_noc_pkt_sent [21] = new();
                  local_noc_pkt_sent [21].header_destination_address  = vLocalToNoC[21].locl__noc__dp_data     ;
                  local_noc_pkt_sent [21].header_source               = 21                                     ;
                  local_noc_pkt_sent [21].header_address_type         = vLocalToNoC[21].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [21].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [21].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 21, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [21]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 22
              @(vLocalToNoC[22].cb_p);
              if ((vLocalToNoC[22].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[22].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 22);
                  local_noc_pkt_sent [22] = new();
                  local_noc_pkt_sent [22].header_destination_address  = vLocalToNoC[22].locl__noc__dp_data     ;
                  local_noc_pkt_sent [22].header_source               = 22                                     ;
                  local_noc_pkt_sent [22].header_address_type         = vLocalToNoC[22].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [22].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [22].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 22, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [22]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 23
              @(vLocalToNoC[23].cb_p);
              if ((vLocalToNoC[23].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[23].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 23);
                  local_noc_pkt_sent [23] = new();
                  local_noc_pkt_sent [23].header_destination_address  = vLocalToNoC[23].locl__noc__dp_data     ;
                  local_noc_pkt_sent [23].header_source               = 23                                     ;
                  local_noc_pkt_sent [23].header_address_type         = vLocalToNoC[23].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [23].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [23].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 23, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [23]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 24
              @(vLocalToNoC[24].cb_p);
              if ((vLocalToNoC[24].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[24].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 24);
                  local_noc_pkt_sent [24] = new();
                  local_noc_pkt_sent [24].header_destination_address  = vLocalToNoC[24].locl__noc__dp_data     ;
                  local_noc_pkt_sent [24].header_source               = 24                                     ;
                  local_noc_pkt_sent [24].header_address_type         = vLocalToNoC[24].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [24].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [24].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 24, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [24]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 25
              @(vLocalToNoC[25].cb_p);
              if ((vLocalToNoC[25].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[25].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 25);
                  local_noc_pkt_sent [25] = new();
                  local_noc_pkt_sent [25].header_destination_address  = vLocalToNoC[25].locl__noc__dp_data     ;
                  local_noc_pkt_sent [25].header_source               = 25                                     ;
                  local_noc_pkt_sent [25].header_address_type         = vLocalToNoC[25].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [25].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [25].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 25, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [25]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 26
              @(vLocalToNoC[26].cb_p);
              if ((vLocalToNoC[26].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[26].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 26);
                  local_noc_pkt_sent [26] = new();
                  local_noc_pkt_sent [26].header_destination_address  = vLocalToNoC[26].locl__noc__dp_data     ;
                  local_noc_pkt_sent [26].header_source               = 26                                     ;
                  local_noc_pkt_sent [26].header_address_type         = vLocalToNoC[26].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [26].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [26].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 26, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [26]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 27
              @(vLocalToNoC[27].cb_p);
              if ((vLocalToNoC[27].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[27].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 27);
                  local_noc_pkt_sent [27] = new();
                  local_noc_pkt_sent [27].header_destination_address  = vLocalToNoC[27].locl__noc__dp_data     ;
                  local_noc_pkt_sent [27].header_source               = 27                                     ;
                  local_noc_pkt_sent [27].header_address_type         = vLocalToNoC[27].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [27].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [27].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 27, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [27]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 28
              @(vLocalToNoC[28].cb_p);
              if ((vLocalToNoC[28].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[28].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 28);
                  local_noc_pkt_sent [28] = new();
                  local_noc_pkt_sent [28].header_destination_address  = vLocalToNoC[28].locl__noc__dp_data     ;
                  local_noc_pkt_sent [28].header_source               = 28                                     ;
                  local_noc_pkt_sent [28].header_address_type         = vLocalToNoC[28].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [28].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [28].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 28, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [28]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 29
              @(vLocalToNoC[29].cb_p);
              if ((vLocalToNoC[29].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[29].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 29);
                  local_noc_pkt_sent [29] = new();
                  local_noc_pkt_sent [29].header_destination_address  = vLocalToNoC[29].locl__noc__dp_data     ;
                  local_noc_pkt_sent [29].header_source               = 29                                     ;
                  local_noc_pkt_sent [29].header_address_type         = vLocalToNoC[29].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [29].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [29].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 29, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [29]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 30
              @(vLocalToNoC[30].cb_p);
              if ((vLocalToNoC[30].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[30].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 30);
                  local_noc_pkt_sent [30] = new();
                  local_noc_pkt_sent [30].header_destination_address  = vLocalToNoC[30].locl__noc__dp_data     ;
                  local_noc_pkt_sent [30].header_source               = 30                                     ;
                  local_noc_pkt_sent [30].header_address_type         = vLocalToNoC[30].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [30].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [30].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 30, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [30]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 31
              @(vLocalToNoC[31].cb_p);
              if ((vLocalToNoC[31].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[31].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 31);
                  local_noc_pkt_sent [31] = new();
                  local_noc_pkt_sent [31].header_destination_address  = vLocalToNoC[31].locl__noc__dp_data     ;
                  local_noc_pkt_sent [31].header_source               = 31                                     ;
                  local_noc_pkt_sent [31].header_address_type         = vLocalToNoC[31].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [31].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [31].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 31, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [31]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 32
              @(vLocalToNoC[32].cb_p);
              if ((vLocalToNoC[32].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[32].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 32);
                  local_noc_pkt_sent [32] = new();
                  local_noc_pkt_sent [32].header_destination_address  = vLocalToNoC[32].locl__noc__dp_data     ;
                  local_noc_pkt_sent [32].header_source               = 32                                     ;
                  local_noc_pkt_sent [32].header_address_type         = vLocalToNoC[32].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [32].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [32].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 32, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [32]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 33
              @(vLocalToNoC[33].cb_p);
              if ((vLocalToNoC[33].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[33].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 33);
                  local_noc_pkt_sent [33] = new();
                  local_noc_pkt_sent [33].header_destination_address  = vLocalToNoC[33].locl__noc__dp_data     ;
                  local_noc_pkt_sent [33].header_source               = 33                                     ;
                  local_noc_pkt_sent [33].header_address_type         = vLocalToNoC[33].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [33].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [33].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 33, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [33]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 34
              @(vLocalToNoC[34].cb_p);
              if ((vLocalToNoC[34].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[34].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 34);
                  local_noc_pkt_sent [34] = new();
                  local_noc_pkt_sent [34].header_destination_address  = vLocalToNoC[34].locl__noc__dp_data     ;
                  local_noc_pkt_sent [34].header_source               = 34                                     ;
                  local_noc_pkt_sent [34].header_address_type         = vLocalToNoC[34].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [34].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [34].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 34, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [34]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 35
              @(vLocalToNoC[35].cb_p);
              if ((vLocalToNoC[35].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[35].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 35);
                  local_noc_pkt_sent [35] = new();
                  local_noc_pkt_sent [35].header_destination_address  = vLocalToNoC[35].locl__noc__dp_data     ;
                  local_noc_pkt_sent [35].header_source               = 35                                     ;
                  local_noc_pkt_sent [35].header_address_type         = vLocalToNoC[35].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [35].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [35].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 35, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [35]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 36
              @(vLocalToNoC[36].cb_p);
              if ((vLocalToNoC[36].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[36].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 36);
                  local_noc_pkt_sent [36] = new();
                  local_noc_pkt_sent [36].header_destination_address  = vLocalToNoC[36].locl__noc__dp_data     ;
                  local_noc_pkt_sent [36].header_source               = 36                                     ;
                  local_noc_pkt_sent [36].header_address_type         = vLocalToNoC[36].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [36].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [36].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 36, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [36]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 37
              @(vLocalToNoC[37].cb_p);
              if ((vLocalToNoC[37].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[37].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 37);
                  local_noc_pkt_sent [37] = new();
                  local_noc_pkt_sent [37].header_destination_address  = vLocalToNoC[37].locl__noc__dp_data     ;
                  local_noc_pkt_sent [37].header_source               = 37                                     ;
                  local_noc_pkt_sent [37].header_address_type         = vLocalToNoC[37].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [37].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [37].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 37, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [37]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 38
              @(vLocalToNoC[38].cb_p);
              if ((vLocalToNoC[38].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[38].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 38);
                  local_noc_pkt_sent [38] = new();
                  local_noc_pkt_sent [38].header_destination_address  = vLocalToNoC[38].locl__noc__dp_data     ;
                  local_noc_pkt_sent [38].header_source               = 38                                     ;
                  local_noc_pkt_sent [38].header_address_type         = vLocalToNoC[38].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [38].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [38].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 38, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [38]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 39
              @(vLocalToNoC[39].cb_p);
              if ((vLocalToNoC[39].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[39].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 39);
                  local_noc_pkt_sent [39] = new();
                  local_noc_pkt_sent [39].header_destination_address  = vLocalToNoC[39].locl__noc__dp_data     ;
                  local_noc_pkt_sent [39].header_source               = 39                                     ;
                  local_noc_pkt_sent [39].header_address_type         = vLocalToNoC[39].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [39].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [39].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 39, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [39]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 40
              @(vLocalToNoC[40].cb_p);
              if ((vLocalToNoC[40].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[40].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 40);
                  local_noc_pkt_sent [40] = new();
                  local_noc_pkt_sent [40].header_destination_address  = vLocalToNoC[40].locl__noc__dp_data     ;
                  local_noc_pkt_sent [40].header_source               = 40                                     ;
                  local_noc_pkt_sent [40].header_address_type         = vLocalToNoC[40].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [40].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [40].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 40, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [40]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 41
              @(vLocalToNoC[41].cb_p);
              if ((vLocalToNoC[41].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[41].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 41);
                  local_noc_pkt_sent [41] = new();
                  local_noc_pkt_sent [41].header_destination_address  = vLocalToNoC[41].locl__noc__dp_data     ;
                  local_noc_pkt_sent [41].header_source               = 41                                     ;
                  local_noc_pkt_sent [41].header_address_type         = vLocalToNoC[41].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [41].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [41].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 41, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [41]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 42
              @(vLocalToNoC[42].cb_p);
              if ((vLocalToNoC[42].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[42].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 42);
                  local_noc_pkt_sent [42] = new();
                  local_noc_pkt_sent [42].header_destination_address  = vLocalToNoC[42].locl__noc__dp_data     ;
                  local_noc_pkt_sent [42].header_source               = 42                                     ;
                  local_noc_pkt_sent [42].header_address_type         = vLocalToNoC[42].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [42].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [42].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 42, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [42]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 43
              @(vLocalToNoC[43].cb_p);
              if ((vLocalToNoC[43].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[43].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 43);
                  local_noc_pkt_sent [43] = new();
                  local_noc_pkt_sent [43].header_destination_address  = vLocalToNoC[43].locl__noc__dp_data     ;
                  local_noc_pkt_sent [43].header_source               = 43                                     ;
                  local_noc_pkt_sent [43].header_address_type         = vLocalToNoC[43].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [43].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [43].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 43, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [43]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 44
              @(vLocalToNoC[44].cb_p);
              if ((vLocalToNoC[44].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[44].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 44);
                  local_noc_pkt_sent [44] = new();
                  local_noc_pkt_sent [44].header_destination_address  = vLocalToNoC[44].locl__noc__dp_data     ;
                  local_noc_pkt_sent [44].header_source               = 44                                     ;
                  local_noc_pkt_sent [44].header_address_type         = vLocalToNoC[44].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [44].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [44].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 44, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [44]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 45
              @(vLocalToNoC[45].cb_p);
              if ((vLocalToNoC[45].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[45].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 45);
                  local_noc_pkt_sent [45] = new();
                  local_noc_pkt_sent [45].header_destination_address  = vLocalToNoC[45].locl__noc__dp_data     ;
                  local_noc_pkt_sent [45].header_source               = 45                                     ;
                  local_noc_pkt_sent [45].header_address_type         = vLocalToNoC[45].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [45].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [45].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 45, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [45]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 46
              @(vLocalToNoC[46].cb_p);
              if ((vLocalToNoC[46].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[46].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 46);
                  local_noc_pkt_sent [46] = new();
                  local_noc_pkt_sent [46].header_destination_address  = vLocalToNoC[46].locl__noc__dp_data     ;
                  local_noc_pkt_sent [46].header_source               = 46                                     ;
                  local_noc_pkt_sent [46].header_address_type         = vLocalToNoC[46].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [46].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [46].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 46, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [46]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 47
              @(vLocalToNoC[47].cb_p);
              if ((vLocalToNoC[47].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[47].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 47);
                  local_noc_pkt_sent [47] = new();
                  local_noc_pkt_sent [47].header_destination_address  = vLocalToNoC[47].locl__noc__dp_data     ;
                  local_noc_pkt_sent [47].header_source               = 47                                     ;
                  local_noc_pkt_sent [47].header_address_type         = vLocalToNoC[47].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [47].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [47].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 47, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [47]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 48
              @(vLocalToNoC[48].cb_p);
              if ((vLocalToNoC[48].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[48].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 48);
                  local_noc_pkt_sent [48] = new();
                  local_noc_pkt_sent [48].header_destination_address  = vLocalToNoC[48].locl__noc__dp_data     ;
                  local_noc_pkt_sent [48].header_source               = 48                                     ;
                  local_noc_pkt_sent [48].header_address_type         = vLocalToNoC[48].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [48].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [48].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 48, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [48]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 49
              @(vLocalToNoC[49].cb_p);
              if ((vLocalToNoC[49].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[49].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 49);
                  local_noc_pkt_sent [49] = new();
                  local_noc_pkt_sent [49].header_destination_address  = vLocalToNoC[49].locl__noc__dp_data     ;
                  local_noc_pkt_sent [49].header_source               = 49                                     ;
                  local_noc_pkt_sent [49].header_address_type         = vLocalToNoC[49].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [49].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [49].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 49, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [49]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 50
              @(vLocalToNoC[50].cb_p);
              if ((vLocalToNoC[50].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[50].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 50);
                  local_noc_pkt_sent [50] = new();
                  local_noc_pkt_sent [50].header_destination_address  = vLocalToNoC[50].locl__noc__dp_data     ;
                  local_noc_pkt_sent [50].header_source               = 50                                     ;
                  local_noc_pkt_sent [50].header_address_type         = vLocalToNoC[50].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [50].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [50].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 50, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [50]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 51
              @(vLocalToNoC[51].cb_p);
              if ((vLocalToNoC[51].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[51].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 51);
                  local_noc_pkt_sent [51] = new();
                  local_noc_pkt_sent [51].header_destination_address  = vLocalToNoC[51].locl__noc__dp_data     ;
                  local_noc_pkt_sent [51].header_source               = 51                                     ;
                  local_noc_pkt_sent [51].header_address_type         = vLocalToNoC[51].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [51].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [51].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 51, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [51]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 52
              @(vLocalToNoC[52].cb_p);
              if ((vLocalToNoC[52].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[52].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 52);
                  local_noc_pkt_sent [52] = new();
                  local_noc_pkt_sent [52].header_destination_address  = vLocalToNoC[52].locl__noc__dp_data     ;
                  local_noc_pkt_sent [52].header_source               = 52                                     ;
                  local_noc_pkt_sent [52].header_address_type         = vLocalToNoC[52].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [52].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [52].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 52, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [52]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 53
              @(vLocalToNoC[53].cb_p);
              if ((vLocalToNoC[53].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[53].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 53);
                  local_noc_pkt_sent [53] = new();
                  local_noc_pkt_sent [53].header_destination_address  = vLocalToNoC[53].locl__noc__dp_data     ;
                  local_noc_pkt_sent [53].header_source               = 53                                     ;
                  local_noc_pkt_sent [53].header_address_type         = vLocalToNoC[53].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [53].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [53].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 53, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [53]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 54
              @(vLocalToNoC[54].cb_p);
              if ((vLocalToNoC[54].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[54].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 54);
                  local_noc_pkt_sent [54] = new();
                  local_noc_pkt_sent [54].header_destination_address  = vLocalToNoC[54].locl__noc__dp_data     ;
                  local_noc_pkt_sent [54].header_source               = 54                                     ;
                  local_noc_pkt_sent [54].header_address_type         = vLocalToNoC[54].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [54].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [54].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 54, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [54]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 55
              @(vLocalToNoC[55].cb_p);
              if ((vLocalToNoC[55].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[55].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 55);
                  local_noc_pkt_sent [55] = new();
                  local_noc_pkt_sent [55].header_destination_address  = vLocalToNoC[55].locl__noc__dp_data     ;
                  local_noc_pkt_sent [55].header_source               = 55                                     ;
                  local_noc_pkt_sent [55].header_address_type         = vLocalToNoC[55].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [55].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [55].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 55, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [55]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 56
              @(vLocalToNoC[56].cb_p);
              if ((vLocalToNoC[56].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[56].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 56);
                  local_noc_pkt_sent [56] = new();
                  local_noc_pkt_sent [56].header_destination_address  = vLocalToNoC[56].locl__noc__dp_data     ;
                  local_noc_pkt_sent [56].header_source               = 56                                     ;
                  local_noc_pkt_sent [56].header_address_type         = vLocalToNoC[56].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [56].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [56].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 56, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [56]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 57
              @(vLocalToNoC[57].cb_p);
              if ((vLocalToNoC[57].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[57].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 57);
                  local_noc_pkt_sent [57] = new();
                  local_noc_pkt_sent [57].header_destination_address  = vLocalToNoC[57].locl__noc__dp_data     ;
                  local_noc_pkt_sent [57].header_source               = 57                                     ;
                  local_noc_pkt_sent [57].header_address_type         = vLocalToNoC[57].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [57].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [57].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 57, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [57]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 58
              @(vLocalToNoC[58].cb_p);
              if ((vLocalToNoC[58].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[58].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 58);
                  local_noc_pkt_sent [58] = new();
                  local_noc_pkt_sent [58].header_destination_address  = vLocalToNoC[58].locl__noc__dp_data     ;
                  local_noc_pkt_sent [58].header_source               = 58                                     ;
                  local_noc_pkt_sent [58].header_address_type         = vLocalToNoC[58].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [58].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [58].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 58, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [58]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 59
              @(vLocalToNoC[59].cb_p);
              if ((vLocalToNoC[59].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[59].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 59);
                  local_noc_pkt_sent [59] = new();
                  local_noc_pkt_sent [59].header_destination_address  = vLocalToNoC[59].locl__noc__dp_data     ;
                  local_noc_pkt_sent [59].header_source               = 59                                     ;
                  local_noc_pkt_sent [59].header_address_type         = vLocalToNoC[59].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [59].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [59].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 59, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [59]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 60
              @(vLocalToNoC[60].cb_p);
              if ((vLocalToNoC[60].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[60].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 60);
                  local_noc_pkt_sent [60] = new();
                  local_noc_pkt_sent [60].header_destination_address  = vLocalToNoC[60].locl__noc__dp_data     ;
                  local_noc_pkt_sent [60].header_source               = 60                                     ;
                  local_noc_pkt_sent [60].header_address_type         = vLocalToNoC[60].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [60].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [60].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 60, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [60]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 61
              @(vLocalToNoC[61].cb_p);
              if ((vLocalToNoC[61].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[61].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 61);
                  local_noc_pkt_sent [61] = new();
                  local_noc_pkt_sent [61].header_destination_address  = vLocalToNoC[61].locl__noc__dp_data     ;
                  local_noc_pkt_sent [61].header_source               = 61                                     ;
                  local_noc_pkt_sent [61].header_address_type         = vLocalToNoC[61].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [61].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [61].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 61, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [61]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 62
              @(vLocalToNoC[62].cb_p);
              if ((vLocalToNoC[62].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[62].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 62);
                  local_noc_pkt_sent [62] = new();
                  local_noc_pkt_sent [62].header_destination_address  = vLocalToNoC[62].locl__noc__dp_data     ;
                  local_noc_pkt_sent [62].header_source               = 62                                     ;
                  local_noc_pkt_sent [62].header_address_type         = vLocalToNoC[62].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [62].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [62].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 62, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [62]);
                        end
                    end
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets sent from manager 63
              @(vLocalToNoC[63].cb_p);
              if ((vLocalToNoC[63].locl__noc__dp_valid == 1'b1) && (vLocalToNoC[63].locl__noc__dp_cntl == 2'b01))
                begin
                  //$display ("@%0t::%s:%0d:: INFO: Packet being sent from {%0d}", $time, `__FILE__, `__LINE__, 63);
                  local_noc_pkt_sent [63] = new();
                  local_noc_pkt_sent [63].header_destination_address  = vLocalToNoC[63].locl__noc__dp_data     ;
                  local_noc_pkt_sent [63].header_source               = 63                                     ;
                  local_noc_pkt_sent [63].header_address_type         = vLocalToNoC[63].locl__noc__dp_desttype ;
                  local_noc_pkt_sent [63].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  // determine all destination and place packet in their mailbox
                  for (int dm=0; dm<`MGR_ARRAY_NUM_OF_MGR; dm++) 
                    begin
                      if (local_noc_pkt_sent [63].header_destination_address[dm] == 1'b1)
                        begin
                          $display ("@%0t::%s:%0d:: INFO: Packet sent from {%0d} to {%0d}", $time, `__FILE__, `__LINE__, 63, dm);
                          mgr2noc_p [dm].put(local_noc_pkt_sent [63]);
                        end
                    end
                end
            end
        end
    