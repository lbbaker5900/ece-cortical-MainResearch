
  assign   pe0__stu__valid                =  pe_inst[0].pe__stu__valid     ;
  assign   pe0__stu__cntl                 =  pe_inst[0].pe__stu__cntl      ;
  assign   pe_inst[0].stu__pe__ready      =  stu__pe0__ready               ;
  assign   pe0__stu__type                 =  pe_inst[0].pe__stu__type      ;
  assign   pe0__stu__data                 =  pe_inst[0].pe__stu__data      ;
  assign   pe0__stu__oob_data             =  pe_inst[0].pe__stu__oob_data  ;

  assign   pe1__stu__valid                =  pe_inst[1].pe__stu__valid     ;
  assign   pe1__stu__cntl                 =  pe_inst[1].pe__stu__cntl      ;
  assign   pe_inst[1].stu__pe__ready      =  stu__pe1__ready               ;
  assign   pe1__stu__type                 =  pe_inst[1].pe__stu__type      ;
  assign   pe1__stu__data                 =  pe_inst[1].pe__stu__data      ;
  assign   pe1__stu__oob_data             =  pe_inst[1].pe__stu__oob_data  ;

  assign   pe2__stu__valid                =  pe_inst[2].pe__stu__valid     ;
  assign   pe2__stu__cntl                 =  pe_inst[2].pe__stu__cntl      ;
  assign   pe_inst[2].stu__pe__ready      =  stu__pe2__ready               ;
  assign   pe2__stu__type                 =  pe_inst[2].pe__stu__type      ;
  assign   pe2__stu__data                 =  pe_inst[2].pe__stu__data      ;
  assign   pe2__stu__oob_data             =  pe_inst[2].pe__stu__oob_data  ;

  assign   pe3__stu__valid                =  pe_inst[3].pe__stu__valid     ;
  assign   pe3__stu__cntl                 =  pe_inst[3].pe__stu__cntl      ;
  assign   pe_inst[3].stu__pe__ready      =  stu__pe3__ready               ;
  assign   pe3__stu__type                 =  pe_inst[3].pe__stu__type      ;
  assign   pe3__stu__data                 =  pe_inst[3].pe__stu__data      ;
  assign   pe3__stu__oob_data             =  pe_inst[3].pe__stu__oob_data  ;

