
//------------------------------------------------
// MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_LOCAL_INPUT_QUEUE_CONTROL_STATE width
//------------------------------------------------
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_STATE_MSB            10
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_STATE_LSB            0
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_STATE_SIZE           (`MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_STATE_MSB - `MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_STATE_LSB +1)
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_STATE_RANGE           `MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_STATE_MSB : `MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_STATE_LSB

//------------------------------------------------------------------------------------------------
//------------------------------------------------
// MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL state machine states
//------------------------------------------------

`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_WAIT        11'd1
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_TRANSFER_LOCAL  11'd2
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_ACK_LOCAL   11'd4
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_TRANSFER_PORT0  11'd8
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_ACK_PORT0   11'd16
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_TRANSFER_PORT1  11'd32
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_ACK_PORT1   11'd64
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_TRANSFER_PORT2  11'd128
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_ACK_PORT2   11'd256
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_TRANSFER_PORT3  11'd512
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_ACK_PORT3   11'd1024