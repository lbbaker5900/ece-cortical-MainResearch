
    assign reg__sdp__lane0_ready    =  reg__scntl__lane0_ready  ;
    assign scntl__reg__lane0_valid  =  sdp__reg__lane0_valid    ;
    assign scntl__reg__lane0_data   =  sdp__reg__lane0_data     ;

    assign reg__sdp__lane1_ready    =  reg__scntl__lane1_ready  ;
    assign scntl__reg__lane1_valid  =  sdp__reg__lane1_valid    ;
    assign scntl__reg__lane1_data   =  sdp__reg__lane1_data     ;

    assign reg__sdp__lane2_ready    =  reg__scntl__lane2_ready  ;
    assign scntl__reg__lane2_valid  =  sdp__reg__lane2_valid    ;
    assign scntl__reg__lane2_data   =  sdp__reg__lane2_data     ;

    assign reg__sdp__lane3_ready    =  reg__scntl__lane3_ready  ;
    assign scntl__reg__lane3_valid  =  sdp__reg__lane3_valid    ;
    assign scntl__reg__lane3_data   =  sdp__reg__lane3_data     ;

    assign reg__sdp__lane4_ready    =  reg__scntl__lane4_ready  ;
    assign scntl__reg__lane4_valid  =  sdp__reg__lane4_valid    ;
    assign scntl__reg__lane4_data   =  sdp__reg__lane4_data     ;

    assign reg__sdp__lane5_ready    =  reg__scntl__lane5_ready  ;
    assign scntl__reg__lane5_valid  =  sdp__reg__lane5_valid    ;
    assign scntl__reg__lane5_data   =  sdp__reg__lane5_data     ;

    assign reg__sdp__lane6_ready    =  reg__scntl__lane6_ready  ;
    assign scntl__reg__lane6_valid  =  sdp__reg__lane6_valid    ;
    assign scntl__reg__lane6_data   =  sdp__reg__lane6_data     ;

    assign reg__sdp__lane7_ready    =  reg__scntl__lane7_ready  ;
    assign scntl__reg__lane7_valid  =  sdp__reg__lane7_valid    ;
    assign scntl__reg__lane7_data   =  sdp__reg__lane7_data     ;

    assign reg__sdp__lane8_ready    =  reg__scntl__lane8_ready  ;
    assign scntl__reg__lane8_valid  =  sdp__reg__lane8_valid    ;
    assign scntl__reg__lane8_data   =  sdp__reg__lane8_data     ;

    assign reg__sdp__lane9_ready    =  reg__scntl__lane9_ready  ;
    assign scntl__reg__lane9_valid  =  sdp__reg__lane9_valid    ;
    assign scntl__reg__lane9_data   =  sdp__reg__lane9_data     ;

    assign reg__sdp__lane10_ready    =  reg__scntl__lane10_ready  ;
    assign scntl__reg__lane10_valid  =  sdp__reg__lane10_valid    ;
    assign scntl__reg__lane10_data   =  sdp__reg__lane10_data     ;

    assign reg__sdp__lane11_ready    =  reg__scntl__lane11_ready  ;
    assign scntl__reg__lane11_valid  =  sdp__reg__lane11_valid    ;
    assign scntl__reg__lane11_data   =  sdp__reg__lane11_data     ;

    assign reg__sdp__lane12_ready    =  reg__scntl__lane12_ready  ;
    assign scntl__reg__lane12_valid  =  sdp__reg__lane12_valid    ;
    assign scntl__reg__lane12_data   =  sdp__reg__lane12_data     ;

    assign reg__sdp__lane13_ready    =  reg__scntl__lane13_ready  ;
    assign scntl__reg__lane13_valid  =  sdp__reg__lane13_valid    ;
    assign scntl__reg__lane13_data   =  sdp__reg__lane13_data     ;

    assign reg__sdp__lane14_ready    =  reg__scntl__lane14_ready  ;
    assign scntl__reg__lane14_valid  =  sdp__reg__lane14_valid    ;
    assign scntl__reg__lane14_data   =  sdp__reg__lane14_data     ;

    assign reg__sdp__lane15_ready    =  reg__scntl__lane15_ready  ;
    assign scntl__reg__lane15_valid  =  sdp__reg__lane15_valid    ;
    assign scntl__reg__lane15_data   =  sdp__reg__lane15_data     ;

    assign reg__sdp__lane16_ready    =  reg__scntl__lane16_ready  ;
    assign scntl__reg__lane16_valid  =  sdp__reg__lane16_valid    ;
    assign scntl__reg__lane16_data   =  sdp__reg__lane16_data     ;

    assign reg__sdp__lane17_ready    =  reg__scntl__lane17_ready  ;
    assign scntl__reg__lane17_valid  =  sdp__reg__lane17_valid    ;
    assign scntl__reg__lane17_data   =  sdp__reg__lane17_data     ;

    assign reg__sdp__lane18_ready    =  reg__scntl__lane18_ready  ;
    assign scntl__reg__lane18_valid  =  sdp__reg__lane18_valid    ;
    assign scntl__reg__lane18_data   =  sdp__reg__lane18_data     ;

    assign reg__sdp__lane19_ready    =  reg__scntl__lane19_ready  ;
    assign scntl__reg__lane19_valid  =  sdp__reg__lane19_valid    ;
    assign scntl__reg__lane19_data   =  sdp__reg__lane19_data     ;

    assign reg__sdp__lane20_ready    =  reg__scntl__lane20_ready  ;
    assign scntl__reg__lane20_valid  =  sdp__reg__lane20_valid    ;
    assign scntl__reg__lane20_data   =  sdp__reg__lane20_data     ;

    assign reg__sdp__lane21_ready    =  reg__scntl__lane21_ready  ;
    assign scntl__reg__lane21_valid  =  sdp__reg__lane21_valid    ;
    assign scntl__reg__lane21_data   =  sdp__reg__lane21_data     ;

    assign reg__sdp__lane22_ready    =  reg__scntl__lane22_ready  ;
    assign scntl__reg__lane22_valid  =  sdp__reg__lane22_valid    ;
    assign scntl__reg__lane22_data   =  sdp__reg__lane22_data     ;

    assign reg__sdp__lane23_ready    =  reg__scntl__lane23_ready  ;
    assign scntl__reg__lane23_valid  =  sdp__reg__lane23_valid    ;
    assign scntl__reg__lane23_data   =  sdp__reg__lane23_data     ;

    assign reg__sdp__lane24_ready    =  reg__scntl__lane24_ready  ;
    assign scntl__reg__lane24_valid  =  sdp__reg__lane24_valid    ;
    assign scntl__reg__lane24_data   =  sdp__reg__lane24_data     ;

    assign reg__sdp__lane25_ready    =  reg__scntl__lane25_ready  ;
    assign scntl__reg__lane25_valid  =  sdp__reg__lane25_valid    ;
    assign scntl__reg__lane25_data   =  sdp__reg__lane25_data     ;

    assign reg__sdp__lane26_ready    =  reg__scntl__lane26_ready  ;
    assign scntl__reg__lane26_valid  =  sdp__reg__lane26_valid    ;
    assign scntl__reg__lane26_data   =  sdp__reg__lane26_data     ;

    assign reg__sdp__lane27_ready    =  reg__scntl__lane27_ready  ;
    assign scntl__reg__lane27_valid  =  sdp__reg__lane27_valid    ;
    assign scntl__reg__lane27_data   =  sdp__reg__lane27_data     ;

    assign reg__sdp__lane28_ready    =  reg__scntl__lane28_ready  ;
    assign scntl__reg__lane28_valid  =  sdp__reg__lane28_valid    ;
    assign scntl__reg__lane28_data   =  sdp__reg__lane28_data     ;

    assign reg__sdp__lane29_ready    =  reg__scntl__lane29_ready  ;
    assign scntl__reg__lane29_valid  =  sdp__reg__lane29_valid    ;
    assign scntl__reg__lane29_data   =  sdp__reg__lane29_data     ;

    assign reg__sdp__lane30_ready    =  reg__scntl__lane30_ready  ;
    assign scntl__reg__lane30_valid  =  sdp__reg__lane30_valid    ;
    assign scntl__reg__lane30_data   =  sdp__reg__lane30_data     ;

    assign reg__sdp__lane31_ready    =  reg__scntl__lane31_ready  ;
    assign scntl__reg__lane31_valid  =  sdp__reg__lane31_valid    ;
    assign scntl__reg__lane31_data   =  sdp__reg__lane31_data     ;

