
        // PE 0, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane0_strm0_ready         ( DownstreamStackBusLane[0][0].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane0_strm0_cntl          ( DownstreamStackBusLane[0][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane0_strm0_data          ( DownstreamStackBusLane[0][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane0_strm0_data_valid    ( DownstreamStackBusLane[0][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane0_strm1_ready         ( DownstreamStackBusLane[0][0].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane0_strm1_cntl          ( DownstreamStackBusLane[0][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane0_strm1_data          ( DownstreamStackBusLane[0][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane0_strm1_data_valid    ( DownstreamStackBusLane[0][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane1_strm0_ready         ( DownstreamStackBusLane[0][1].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane1_strm0_cntl          ( DownstreamStackBusLane[0][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane1_strm0_data          ( DownstreamStackBusLane[0][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane1_strm0_data_valid    ( DownstreamStackBusLane[0][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane1_strm1_ready         ( DownstreamStackBusLane[0][1].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane1_strm1_cntl          ( DownstreamStackBusLane[0][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane1_strm1_data          ( DownstreamStackBusLane[0][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane1_strm1_data_valid    ( DownstreamStackBusLane[0][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane2_strm0_ready         ( DownstreamStackBusLane[0][2].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane2_strm0_cntl          ( DownstreamStackBusLane[0][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane2_strm0_data          ( DownstreamStackBusLane[0][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane2_strm0_data_valid    ( DownstreamStackBusLane[0][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane2_strm1_ready         ( DownstreamStackBusLane[0][2].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane2_strm1_cntl          ( DownstreamStackBusLane[0][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane2_strm1_data          ( DownstreamStackBusLane[0][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane2_strm1_data_valid    ( DownstreamStackBusLane[0][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane3_strm0_ready         ( DownstreamStackBusLane[0][3].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane3_strm0_cntl          ( DownstreamStackBusLane[0][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane3_strm0_data          ( DownstreamStackBusLane[0][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane3_strm0_data_valid    ( DownstreamStackBusLane[0][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane3_strm1_ready         ( DownstreamStackBusLane[0][3].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane3_strm1_cntl          ( DownstreamStackBusLane[0][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane3_strm1_data          ( DownstreamStackBusLane[0][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane3_strm1_data_valid    ( DownstreamStackBusLane[0][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane4_strm0_ready         ( DownstreamStackBusLane[0][4].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane4_strm0_cntl          ( DownstreamStackBusLane[0][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane4_strm0_data          ( DownstreamStackBusLane[0][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane4_strm0_data_valid    ( DownstreamStackBusLane[0][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane4_strm1_ready         ( DownstreamStackBusLane[0][4].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane4_strm1_cntl          ( DownstreamStackBusLane[0][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane4_strm1_data          ( DownstreamStackBusLane[0][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane4_strm1_data_valid    ( DownstreamStackBusLane[0][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane5_strm0_ready         ( DownstreamStackBusLane[0][5].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane5_strm0_cntl          ( DownstreamStackBusLane[0][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane5_strm0_data          ( DownstreamStackBusLane[0][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane5_strm0_data_valid    ( DownstreamStackBusLane[0][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane5_strm1_ready         ( DownstreamStackBusLane[0][5].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane5_strm1_cntl          ( DownstreamStackBusLane[0][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane5_strm1_data          ( DownstreamStackBusLane[0][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane5_strm1_data_valid    ( DownstreamStackBusLane[0][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane6_strm0_ready         ( DownstreamStackBusLane[0][6].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane6_strm0_cntl          ( DownstreamStackBusLane[0][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane6_strm0_data          ( DownstreamStackBusLane[0][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane6_strm0_data_valid    ( DownstreamStackBusLane[0][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane6_strm1_ready         ( DownstreamStackBusLane[0][6].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane6_strm1_cntl          ( DownstreamStackBusLane[0][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane6_strm1_data          ( DownstreamStackBusLane[0][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane6_strm1_data_valid    ( DownstreamStackBusLane[0][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane7_strm0_ready         ( DownstreamStackBusLane[0][7].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane7_strm0_cntl          ( DownstreamStackBusLane[0][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane7_strm0_data          ( DownstreamStackBusLane[0][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane7_strm0_data_valid    ( DownstreamStackBusLane[0][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane7_strm1_ready         ( DownstreamStackBusLane[0][7].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane7_strm1_cntl          ( DownstreamStackBusLane[0][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane7_strm1_data          ( DownstreamStackBusLane[0][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane7_strm1_data_valid    ( DownstreamStackBusLane[0][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane8_strm0_ready         ( DownstreamStackBusLane[0][8].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane8_strm0_cntl          ( DownstreamStackBusLane[0][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane8_strm0_data          ( DownstreamStackBusLane[0][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane8_strm0_data_valid    ( DownstreamStackBusLane[0][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane8_strm1_ready         ( DownstreamStackBusLane[0][8].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane8_strm1_cntl          ( DownstreamStackBusLane[0][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane8_strm1_data          ( DownstreamStackBusLane[0][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane8_strm1_data_valid    ( DownstreamStackBusLane[0][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane9_strm0_ready         ( DownstreamStackBusLane[0][9].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane9_strm0_cntl          ( DownstreamStackBusLane[0][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane9_strm0_data          ( DownstreamStackBusLane[0][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane9_strm0_data_valid    ( DownstreamStackBusLane[0][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane9_strm1_ready         ( DownstreamStackBusLane[0][9].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane9_strm1_cntl          ( DownstreamStackBusLane[0][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane9_strm1_data          ( DownstreamStackBusLane[0][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane9_strm1_data_valid    ( DownstreamStackBusLane[0][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane10_strm0_ready         ( DownstreamStackBusLane[0][10].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane10_strm0_cntl          ( DownstreamStackBusLane[0][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane10_strm0_data          ( DownstreamStackBusLane[0][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane10_strm0_data_valid    ( DownstreamStackBusLane[0][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane10_strm1_ready         ( DownstreamStackBusLane[0][10].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane10_strm1_cntl          ( DownstreamStackBusLane[0][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane10_strm1_data          ( DownstreamStackBusLane[0][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane10_strm1_data_valid    ( DownstreamStackBusLane[0][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane11_strm0_ready         ( DownstreamStackBusLane[0][11].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane11_strm0_cntl          ( DownstreamStackBusLane[0][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane11_strm0_data          ( DownstreamStackBusLane[0][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane11_strm0_data_valid    ( DownstreamStackBusLane[0][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane11_strm1_ready         ( DownstreamStackBusLane[0][11].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane11_strm1_cntl          ( DownstreamStackBusLane[0][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane11_strm1_data          ( DownstreamStackBusLane[0][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane11_strm1_data_valid    ( DownstreamStackBusLane[0][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane12_strm0_ready         ( DownstreamStackBusLane[0][12].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane12_strm0_cntl          ( DownstreamStackBusLane[0][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane12_strm0_data          ( DownstreamStackBusLane[0][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane12_strm0_data_valid    ( DownstreamStackBusLane[0][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane12_strm1_ready         ( DownstreamStackBusLane[0][12].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane12_strm1_cntl          ( DownstreamStackBusLane[0][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane12_strm1_data          ( DownstreamStackBusLane[0][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane12_strm1_data_valid    ( DownstreamStackBusLane[0][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane13_strm0_ready         ( DownstreamStackBusLane[0][13].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane13_strm0_cntl          ( DownstreamStackBusLane[0][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane13_strm0_data          ( DownstreamStackBusLane[0][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane13_strm0_data_valid    ( DownstreamStackBusLane[0][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane13_strm1_ready         ( DownstreamStackBusLane[0][13].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane13_strm1_cntl          ( DownstreamStackBusLane[0][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane13_strm1_data          ( DownstreamStackBusLane[0][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane13_strm1_data_valid    ( DownstreamStackBusLane[0][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane14_strm0_ready         ( DownstreamStackBusLane[0][14].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane14_strm0_cntl          ( DownstreamStackBusLane[0][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane14_strm0_data          ( DownstreamStackBusLane[0][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane14_strm0_data_valid    ( DownstreamStackBusLane[0][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane14_strm1_ready         ( DownstreamStackBusLane[0][14].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane14_strm1_cntl          ( DownstreamStackBusLane[0][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane14_strm1_data          ( DownstreamStackBusLane[0][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane14_strm1_data_valid    ( DownstreamStackBusLane[0][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane15_strm0_ready         ( DownstreamStackBusLane[0][15].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane15_strm0_cntl          ( DownstreamStackBusLane[0][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane15_strm0_data          ( DownstreamStackBusLane[0][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane15_strm0_data_valid    ( DownstreamStackBusLane[0][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane15_strm1_ready         ( DownstreamStackBusLane[0][15].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane15_strm1_cntl          ( DownstreamStackBusLane[0][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane15_strm1_data          ( DownstreamStackBusLane[0][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane15_strm1_data_valid    ( DownstreamStackBusLane[0][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane16_strm0_ready         ( DownstreamStackBusLane[0][16].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane16_strm0_cntl          ( DownstreamStackBusLane[0][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane16_strm0_data          ( DownstreamStackBusLane[0][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane16_strm0_data_valid    ( DownstreamStackBusLane[0][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane16_strm1_ready         ( DownstreamStackBusLane[0][16].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane16_strm1_cntl          ( DownstreamStackBusLane[0][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane16_strm1_data          ( DownstreamStackBusLane[0][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane16_strm1_data_valid    ( DownstreamStackBusLane[0][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane17_strm0_ready         ( DownstreamStackBusLane[0][17].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane17_strm0_cntl          ( DownstreamStackBusLane[0][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane17_strm0_data          ( DownstreamStackBusLane[0][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane17_strm0_data_valid    ( DownstreamStackBusLane[0][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane17_strm1_ready         ( DownstreamStackBusLane[0][17].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane17_strm1_cntl          ( DownstreamStackBusLane[0][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane17_strm1_data          ( DownstreamStackBusLane[0][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane17_strm1_data_valid    ( DownstreamStackBusLane[0][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane18_strm0_ready         ( DownstreamStackBusLane[0][18].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane18_strm0_cntl          ( DownstreamStackBusLane[0][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane18_strm0_data          ( DownstreamStackBusLane[0][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane18_strm0_data_valid    ( DownstreamStackBusLane[0][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane18_strm1_ready         ( DownstreamStackBusLane[0][18].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane18_strm1_cntl          ( DownstreamStackBusLane[0][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane18_strm1_data          ( DownstreamStackBusLane[0][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane18_strm1_data_valid    ( DownstreamStackBusLane[0][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane19_strm0_ready         ( DownstreamStackBusLane[0][19].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane19_strm0_cntl          ( DownstreamStackBusLane[0][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane19_strm0_data          ( DownstreamStackBusLane[0][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane19_strm0_data_valid    ( DownstreamStackBusLane[0][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane19_strm1_ready         ( DownstreamStackBusLane[0][19].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane19_strm1_cntl          ( DownstreamStackBusLane[0][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane19_strm1_data          ( DownstreamStackBusLane[0][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane19_strm1_data_valid    ( DownstreamStackBusLane[0][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane20_strm0_ready         ( DownstreamStackBusLane[0][20].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane20_strm0_cntl          ( DownstreamStackBusLane[0][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane20_strm0_data          ( DownstreamStackBusLane[0][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane20_strm0_data_valid    ( DownstreamStackBusLane[0][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane20_strm1_ready         ( DownstreamStackBusLane[0][20].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane20_strm1_cntl          ( DownstreamStackBusLane[0][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane20_strm1_data          ( DownstreamStackBusLane[0][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane20_strm1_data_valid    ( DownstreamStackBusLane[0][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane21_strm0_ready         ( DownstreamStackBusLane[0][21].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane21_strm0_cntl          ( DownstreamStackBusLane[0][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane21_strm0_data          ( DownstreamStackBusLane[0][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane21_strm0_data_valid    ( DownstreamStackBusLane[0][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane21_strm1_ready         ( DownstreamStackBusLane[0][21].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane21_strm1_cntl          ( DownstreamStackBusLane[0][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane21_strm1_data          ( DownstreamStackBusLane[0][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane21_strm1_data_valid    ( DownstreamStackBusLane[0][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane22_strm0_ready         ( DownstreamStackBusLane[0][22].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane22_strm0_cntl          ( DownstreamStackBusLane[0][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane22_strm0_data          ( DownstreamStackBusLane[0][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane22_strm0_data_valid    ( DownstreamStackBusLane[0][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane22_strm1_ready         ( DownstreamStackBusLane[0][22].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane22_strm1_cntl          ( DownstreamStackBusLane[0][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane22_strm1_data          ( DownstreamStackBusLane[0][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane22_strm1_data_valid    ( DownstreamStackBusLane[0][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane23_strm0_ready         ( DownstreamStackBusLane[0][23].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane23_strm0_cntl          ( DownstreamStackBusLane[0][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane23_strm0_data          ( DownstreamStackBusLane[0][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane23_strm0_data_valid    ( DownstreamStackBusLane[0][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane23_strm1_ready         ( DownstreamStackBusLane[0][23].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane23_strm1_cntl          ( DownstreamStackBusLane[0][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane23_strm1_data          ( DownstreamStackBusLane[0][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane23_strm1_data_valid    ( DownstreamStackBusLane[0][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane24_strm0_ready         ( DownstreamStackBusLane[0][24].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane24_strm0_cntl          ( DownstreamStackBusLane[0][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane24_strm0_data          ( DownstreamStackBusLane[0][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane24_strm0_data_valid    ( DownstreamStackBusLane[0][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane24_strm1_ready         ( DownstreamStackBusLane[0][24].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane24_strm1_cntl          ( DownstreamStackBusLane[0][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane24_strm1_data          ( DownstreamStackBusLane[0][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane24_strm1_data_valid    ( DownstreamStackBusLane[0][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane25_strm0_ready         ( DownstreamStackBusLane[0][25].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane25_strm0_cntl          ( DownstreamStackBusLane[0][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane25_strm0_data          ( DownstreamStackBusLane[0][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane25_strm0_data_valid    ( DownstreamStackBusLane[0][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane25_strm1_ready         ( DownstreamStackBusLane[0][25].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane25_strm1_cntl          ( DownstreamStackBusLane[0][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane25_strm1_data          ( DownstreamStackBusLane[0][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane25_strm1_data_valid    ( DownstreamStackBusLane[0][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane26_strm0_ready         ( DownstreamStackBusLane[0][26].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane26_strm0_cntl          ( DownstreamStackBusLane[0][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane26_strm0_data          ( DownstreamStackBusLane[0][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane26_strm0_data_valid    ( DownstreamStackBusLane[0][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane26_strm1_ready         ( DownstreamStackBusLane[0][26].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane26_strm1_cntl          ( DownstreamStackBusLane[0][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane26_strm1_data          ( DownstreamStackBusLane[0][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane26_strm1_data_valid    ( DownstreamStackBusLane[0][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane27_strm0_ready         ( DownstreamStackBusLane[0][27].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane27_strm0_cntl          ( DownstreamStackBusLane[0][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane27_strm0_data          ( DownstreamStackBusLane[0][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane27_strm0_data_valid    ( DownstreamStackBusLane[0][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane27_strm1_ready         ( DownstreamStackBusLane[0][27].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane27_strm1_cntl          ( DownstreamStackBusLane[0][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane27_strm1_data          ( DownstreamStackBusLane[0][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane27_strm1_data_valid    ( DownstreamStackBusLane[0][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane28_strm0_ready         ( DownstreamStackBusLane[0][28].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane28_strm0_cntl          ( DownstreamStackBusLane[0][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane28_strm0_data          ( DownstreamStackBusLane[0][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane28_strm0_data_valid    ( DownstreamStackBusLane[0][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane28_strm1_ready         ( DownstreamStackBusLane[0][28].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane28_strm1_cntl          ( DownstreamStackBusLane[0][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane28_strm1_data          ( DownstreamStackBusLane[0][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane28_strm1_data_valid    ( DownstreamStackBusLane[0][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane29_strm0_ready         ( DownstreamStackBusLane[0][29].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane29_strm0_cntl          ( DownstreamStackBusLane[0][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane29_strm0_data          ( DownstreamStackBusLane[0][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane29_strm0_data_valid    ( DownstreamStackBusLane[0][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane29_strm1_ready         ( DownstreamStackBusLane[0][29].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane29_strm1_cntl          ( DownstreamStackBusLane[0][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane29_strm1_data          ( DownstreamStackBusLane[0][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane29_strm1_data_valid    ( DownstreamStackBusLane[0][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane30_strm0_ready         ( DownstreamStackBusLane[0][30].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane30_strm0_cntl          ( DownstreamStackBusLane[0][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane30_strm0_data          ( DownstreamStackBusLane[0][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane30_strm0_data_valid    ( DownstreamStackBusLane[0][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane30_strm1_ready         ( DownstreamStackBusLane[0][30].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane30_strm1_cntl          ( DownstreamStackBusLane[0][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane30_strm1_data          ( DownstreamStackBusLane[0][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane30_strm1_data_valid    ( DownstreamStackBusLane[0][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 0, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane31_strm0_ready         ( DownstreamStackBusLane[0][31].pe__std__lane_strm0_ready              ),      
        .std__pe0__lane31_strm0_cntl          ( DownstreamStackBusLane[0][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe0__lane31_strm0_data          ( DownstreamStackBusLane[0][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe0__lane31_strm0_data_valid    ( DownstreamStackBusLane[0][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__std__lane31_strm1_ready         ( DownstreamStackBusLane[0][31].pe__std__lane_strm1_ready              ),      
        .std__pe0__lane31_strm1_cntl          ( DownstreamStackBusLane[0][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe0__lane31_strm1_data          ( DownstreamStackBusLane[0][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe0__lane31_strm1_data_valid    ( DownstreamStackBusLane[0][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane0_strm0_ready         ( DownstreamStackBusLane[1][0].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane0_strm0_cntl          ( DownstreamStackBusLane[1][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane0_strm0_data          ( DownstreamStackBusLane[1][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane0_strm0_data_valid    ( DownstreamStackBusLane[1][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane0_strm1_ready         ( DownstreamStackBusLane[1][0].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane0_strm1_cntl          ( DownstreamStackBusLane[1][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane0_strm1_data          ( DownstreamStackBusLane[1][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane0_strm1_data_valid    ( DownstreamStackBusLane[1][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane1_strm0_ready         ( DownstreamStackBusLane[1][1].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane1_strm0_cntl          ( DownstreamStackBusLane[1][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane1_strm0_data          ( DownstreamStackBusLane[1][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane1_strm0_data_valid    ( DownstreamStackBusLane[1][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane1_strm1_ready         ( DownstreamStackBusLane[1][1].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane1_strm1_cntl          ( DownstreamStackBusLane[1][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane1_strm1_data          ( DownstreamStackBusLane[1][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane1_strm1_data_valid    ( DownstreamStackBusLane[1][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane2_strm0_ready         ( DownstreamStackBusLane[1][2].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane2_strm0_cntl          ( DownstreamStackBusLane[1][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane2_strm0_data          ( DownstreamStackBusLane[1][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane2_strm0_data_valid    ( DownstreamStackBusLane[1][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane2_strm1_ready         ( DownstreamStackBusLane[1][2].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane2_strm1_cntl          ( DownstreamStackBusLane[1][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane2_strm1_data          ( DownstreamStackBusLane[1][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane2_strm1_data_valid    ( DownstreamStackBusLane[1][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane3_strm0_ready         ( DownstreamStackBusLane[1][3].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane3_strm0_cntl          ( DownstreamStackBusLane[1][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane3_strm0_data          ( DownstreamStackBusLane[1][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane3_strm0_data_valid    ( DownstreamStackBusLane[1][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane3_strm1_ready         ( DownstreamStackBusLane[1][3].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane3_strm1_cntl          ( DownstreamStackBusLane[1][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane3_strm1_data          ( DownstreamStackBusLane[1][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane3_strm1_data_valid    ( DownstreamStackBusLane[1][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane4_strm0_ready         ( DownstreamStackBusLane[1][4].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane4_strm0_cntl          ( DownstreamStackBusLane[1][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane4_strm0_data          ( DownstreamStackBusLane[1][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane4_strm0_data_valid    ( DownstreamStackBusLane[1][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane4_strm1_ready         ( DownstreamStackBusLane[1][4].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane4_strm1_cntl          ( DownstreamStackBusLane[1][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane4_strm1_data          ( DownstreamStackBusLane[1][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane4_strm1_data_valid    ( DownstreamStackBusLane[1][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane5_strm0_ready         ( DownstreamStackBusLane[1][5].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane5_strm0_cntl          ( DownstreamStackBusLane[1][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane5_strm0_data          ( DownstreamStackBusLane[1][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane5_strm0_data_valid    ( DownstreamStackBusLane[1][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane5_strm1_ready         ( DownstreamStackBusLane[1][5].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane5_strm1_cntl          ( DownstreamStackBusLane[1][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane5_strm1_data          ( DownstreamStackBusLane[1][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane5_strm1_data_valid    ( DownstreamStackBusLane[1][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane6_strm0_ready         ( DownstreamStackBusLane[1][6].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane6_strm0_cntl          ( DownstreamStackBusLane[1][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane6_strm0_data          ( DownstreamStackBusLane[1][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane6_strm0_data_valid    ( DownstreamStackBusLane[1][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane6_strm1_ready         ( DownstreamStackBusLane[1][6].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane6_strm1_cntl          ( DownstreamStackBusLane[1][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane6_strm1_data          ( DownstreamStackBusLane[1][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane6_strm1_data_valid    ( DownstreamStackBusLane[1][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane7_strm0_ready         ( DownstreamStackBusLane[1][7].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane7_strm0_cntl          ( DownstreamStackBusLane[1][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane7_strm0_data          ( DownstreamStackBusLane[1][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane7_strm0_data_valid    ( DownstreamStackBusLane[1][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane7_strm1_ready         ( DownstreamStackBusLane[1][7].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane7_strm1_cntl          ( DownstreamStackBusLane[1][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane7_strm1_data          ( DownstreamStackBusLane[1][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane7_strm1_data_valid    ( DownstreamStackBusLane[1][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane8_strm0_ready         ( DownstreamStackBusLane[1][8].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane8_strm0_cntl          ( DownstreamStackBusLane[1][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane8_strm0_data          ( DownstreamStackBusLane[1][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane8_strm0_data_valid    ( DownstreamStackBusLane[1][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane8_strm1_ready         ( DownstreamStackBusLane[1][8].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane8_strm1_cntl          ( DownstreamStackBusLane[1][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane8_strm1_data          ( DownstreamStackBusLane[1][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane8_strm1_data_valid    ( DownstreamStackBusLane[1][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane9_strm0_ready         ( DownstreamStackBusLane[1][9].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane9_strm0_cntl          ( DownstreamStackBusLane[1][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane9_strm0_data          ( DownstreamStackBusLane[1][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane9_strm0_data_valid    ( DownstreamStackBusLane[1][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane9_strm1_ready         ( DownstreamStackBusLane[1][9].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane9_strm1_cntl          ( DownstreamStackBusLane[1][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane9_strm1_data          ( DownstreamStackBusLane[1][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane9_strm1_data_valid    ( DownstreamStackBusLane[1][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane10_strm0_ready         ( DownstreamStackBusLane[1][10].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane10_strm0_cntl          ( DownstreamStackBusLane[1][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane10_strm0_data          ( DownstreamStackBusLane[1][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane10_strm0_data_valid    ( DownstreamStackBusLane[1][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane10_strm1_ready         ( DownstreamStackBusLane[1][10].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane10_strm1_cntl          ( DownstreamStackBusLane[1][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane10_strm1_data          ( DownstreamStackBusLane[1][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane10_strm1_data_valid    ( DownstreamStackBusLane[1][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane11_strm0_ready         ( DownstreamStackBusLane[1][11].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane11_strm0_cntl          ( DownstreamStackBusLane[1][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane11_strm0_data          ( DownstreamStackBusLane[1][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane11_strm0_data_valid    ( DownstreamStackBusLane[1][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane11_strm1_ready         ( DownstreamStackBusLane[1][11].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane11_strm1_cntl          ( DownstreamStackBusLane[1][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane11_strm1_data          ( DownstreamStackBusLane[1][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane11_strm1_data_valid    ( DownstreamStackBusLane[1][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane12_strm0_ready         ( DownstreamStackBusLane[1][12].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane12_strm0_cntl          ( DownstreamStackBusLane[1][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane12_strm0_data          ( DownstreamStackBusLane[1][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane12_strm0_data_valid    ( DownstreamStackBusLane[1][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane12_strm1_ready         ( DownstreamStackBusLane[1][12].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane12_strm1_cntl          ( DownstreamStackBusLane[1][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane12_strm1_data          ( DownstreamStackBusLane[1][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane12_strm1_data_valid    ( DownstreamStackBusLane[1][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane13_strm0_ready         ( DownstreamStackBusLane[1][13].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane13_strm0_cntl          ( DownstreamStackBusLane[1][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane13_strm0_data          ( DownstreamStackBusLane[1][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane13_strm0_data_valid    ( DownstreamStackBusLane[1][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane13_strm1_ready         ( DownstreamStackBusLane[1][13].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane13_strm1_cntl          ( DownstreamStackBusLane[1][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane13_strm1_data          ( DownstreamStackBusLane[1][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane13_strm1_data_valid    ( DownstreamStackBusLane[1][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane14_strm0_ready         ( DownstreamStackBusLane[1][14].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane14_strm0_cntl          ( DownstreamStackBusLane[1][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane14_strm0_data          ( DownstreamStackBusLane[1][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane14_strm0_data_valid    ( DownstreamStackBusLane[1][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane14_strm1_ready         ( DownstreamStackBusLane[1][14].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane14_strm1_cntl          ( DownstreamStackBusLane[1][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane14_strm1_data          ( DownstreamStackBusLane[1][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane14_strm1_data_valid    ( DownstreamStackBusLane[1][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane15_strm0_ready         ( DownstreamStackBusLane[1][15].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane15_strm0_cntl          ( DownstreamStackBusLane[1][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane15_strm0_data          ( DownstreamStackBusLane[1][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane15_strm0_data_valid    ( DownstreamStackBusLane[1][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane15_strm1_ready         ( DownstreamStackBusLane[1][15].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane15_strm1_cntl          ( DownstreamStackBusLane[1][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane15_strm1_data          ( DownstreamStackBusLane[1][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane15_strm1_data_valid    ( DownstreamStackBusLane[1][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane16_strm0_ready         ( DownstreamStackBusLane[1][16].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane16_strm0_cntl          ( DownstreamStackBusLane[1][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane16_strm0_data          ( DownstreamStackBusLane[1][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane16_strm0_data_valid    ( DownstreamStackBusLane[1][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane16_strm1_ready         ( DownstreamStackBusLane[1][16].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane16_strm1_cntl          ( DownstreamStackBusLane[1][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane16_strm1_data          ( DownstreamStackBusLane[1][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane16_strm1_data_valid    ( DownstreamStackBusLane[1][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane17_strm0_ready         ( DownstreamStackBusLane[1][17].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane17_strm0_cntl          ( DownstreamStackBusLane[1][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane17_strm0_data          ( DownstreamStackBusLane[1][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane17_strm0_data_valid    ( DownstreamStackBusLane[1][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane17_strm1_ready         ( DownstreamStackBusLane[1][17].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane17_strm1_cntl          ( DownstreamStackBusLane[1][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane17_strm1_data          ( DownstreamStackBusLane[1][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane17_strm1_data_valid    ( DownstreamStackBusLane[1][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane18_strm0_ready         ( DownstreamStackBusLane[1][18].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane18_strm0_cntl          ( DownstreamStackBusLane[1][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane18_strm0_data          ( DownstreamStackBusLane[1][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane18_strm0_data_valid    ( DownstreamStackBusLane[1][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane18_strm1_ready         ( DownstreamStackBusLane[1][18].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane18_strm1_cntl          ( DownstreamStackBusLane[1][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane18_strm1_data          ( DownstreamStackBusLane[1][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane18_strm1_data_valid    ( DownstreamStackBusLane[1][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane19_strm0_ready         ( DownstreamStackBusLane[1][19].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane19_strm0_cntl          ( DownstreamStackBusLane[1][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane19_strm0_data          ( DownstreamStackBusLane[1][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane19_strm0_data_valid    ( DownstreamStackBusLane[1][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane19_strm1_ready         ( DownstreamStackBusLane[1][19].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane19_strm1_cntl          ( DownstreamStackBusLane[1][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane19_strm1_data          ( DownstreamStackBusLane[1][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane19_strm1_data_valid    ( DownstreamStackBusLane[1][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane20_strm0_ready         ( DownstreamStackBusLane[1][20].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane20_strm0_cntl          ( DownstreamStackBusLane[1][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane20_strm0_data          ( DownstreamStackBusLane[1][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane20_strm0_data_valid    ( DownstreamStackBusLane[1][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane20_strm1_ready         ( DownstreamStackBusLane[1][20].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane20_strm1_cntl          ( DownstreamStackBusLane[1][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane20_strm1_data          ( DownstreamStackBusLane[1][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane20_strm1_data_valid    ( DownstreamStackBusLane[1][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane21_strm0_ready         ( DownstreamStackBusLane[1][21].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane21_strm0_cntl          ( DownstreamStackBusLane[1][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane21_strm0_data          ( DownstreamStackBusLane[1][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane21_strm0_data_valid    ( DownstreamStackBusLane[1][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane21_strm1_ready         ( DownstreamStackBusLane[1][21].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane21_strm1_cntl          ( DownstreamStackBusLane[1][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane21_strm1_data          ( DownstreamStackBusLane[1][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane21_strm1_data_valid    ( DownstreamStackBusLane[1][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane22_strm0_ready         ( DownstreamStackBusLane[1][22].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane22_strm0_cntl          ( DownstreamStackBusLane[1][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane22_strm0_data          ( DownstreamStackBusLane[1][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane22_strm0_data_valid    ( DownstreamStackBusLane[1][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane22_strm1_ready         ( DownstreamStackBusLane[1][22].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane22_strm1_cntl          ( DownstreamStackBusLane[1][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane22_strm1_data          ( DownstreamStackBusLane[1][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane22_strm1_data_valid    ( DownstreamStackBusLane[1][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane23_strm0_ready         ( DownstreamStackBusLane[1][23].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane23_strm0_cntl          ( DownstreamStackBusLane[1][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane23_strm0_data          ( DownstreamStackBusLane[1][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane23_strm0_data_valid    ( DownstreamStackBusLane[1][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane23_strm1_ready         ( DownstreamStackBusLane[1][23].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane23_strm1_cntl          ( DownstreamStackBusLane[1][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane23_strm1_data          ( DownstreamStackBusLane[1][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane23_strm1_data_valid    ( DownstreamStackBusLane[1][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane24_strm0_ready         ( DownstreamStackBusLane[1][24].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane24_strm0_cntl          ( DownstreamStackBusLane[1][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane24_strm0_data          ( DownstreamStackBusLane[1][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane24_strm0_data_valid    ( DownstreamStackBusLane[1][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane24_strm1_ready         ( DownstreamStackBusLane[1][24].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane24_strm1_cntl          ( DownstreamStackBusLane[1][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane24_strm1_data          ( DownstreamStackBusLane[1][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane24_strm1_data_valid    ( DownstreamStackBusLane[1][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane25_strm0_ready         ( DownstreamStackBusLane[1][25].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane25_strm0_cntl          ( DownstreamStackBusLane[1][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane25_strm0_data          ( DownstreamStackBusLane[1][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane25_strm0_data_valid    ( DownstreamStackBusLane[1][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane25_strm1_ready         ( DownstreamStackBusLane[1][25].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane25_strm1_cntl          ( DownstreamStackBusLane[1][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane25_strm1_data          ( DownstreamStackBusLane[1][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane25_strm1_data_valid    ( DownstreamStackBusLane[1][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane26_strm0_ready         ( DownstreamStackBusLane[1][26].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane26_strm0_cntl          ( DownstreamStackBusLane[1][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane26_strm0_data          ( DownstreamStackBusLane[1][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane26_strm0_data_valid    ( DownstreamStackBusLane[1][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane26_strm1_ready         ( DownstreamStackBusLane[1][26].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane26_strm1_cntl          ( DownstreamStackBusLane[1][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane26_strm1_data          ( DownstreamStackBusLane[1][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane26_strm1_data_valid    ( DownstreamStackBusLane[1][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane27_strm0_ready         ( DownstreamStackBusLane[1][27].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane27_strm0_cntl          ( DownstreamStackBusLane[1][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane27_strm0_data          ( DownstreamStackBusLane[1][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane27_strm0_data_valid    ( DownstreamStackBusLane[1][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane27_strm1_ready         ( DownstreamStackBusLane[1][27].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane27_strm1_cntl          ( DownstreamStackBusLane[1][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane27_strm1_data          ( DownstreamStackBusLane[1][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane27_strm1_data_valid    ( DownstreamStackBusLane[1][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane28_strm0_ready         ( DownstreamStackBusLane[1][28].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane28_strm0_cntl          ( DownstreamStackBusLane[1][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane28_strm0_data          ( DownstreamStackBusLane[1][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane28_strm0_data_valid    ( DownstreamStackBusLane[1][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane28_strm1_ready         ( DownstreamStackBusLane[1][28].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane28_strm1_cntl          ( DownstreamStackBusLane[1][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane28_strm1_data          ( DownstreamStackBusLane[1][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane28_strm1_data_valid    ( DownstreamStackBusLane[1][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane29_strm0_ready         ( DownstreamStackBusLane[1][29].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane29_strm0_cntl          ( DownstreamStackBusLane[1][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane29_strm0_data          ( DownstreamStackBusLane[1][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane29_strm0_data_valid    ( DownstreamStackBusLane[1][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane29_strm1_ready         ( DownstreamStackBusLane[1][29].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane29_strm1_cntl          ( DownstreamStackBusLane[1][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane29_strm1_data          ( DownstreamStackBusLane[1][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane29_strm1_data_valid    ( DownstreamStackBusLane[1][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane30_strm0_ready         ( DownstreamStackBusLane[1][30].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane30_strm0_cntl          ( DownstreamStackBusLane[1][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane30_strm0_data          ( DownstreamStackBusLane[1][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane30_strm0_data_valid    ( DownstreamStackBusLane[1][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane30_strm1_ready         ( DownstreamStackBusLane[1][30].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane30_strm1_cntl          ( DownstreamStackBusLane[1][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane30_strm1_data          ( DownstreamStackBusLane[1][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane30_strm1_data_valid    ( DownstreamStackBusLane[1][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 1, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane31_strm0_ready         ( DownstreamStackBusLane[1][31].pe__std__lane_strm0_ready              ),      
        .std__pe1__lane31_strm0_cntl          ( DownstreamStackBusLane[1][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe1__lane31_strm0_data          ( DownstreamStackBusLane[1][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe1__lane31_strm0_data_valid    ( DownstreamStackBusLane[1][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__std__lane31_strm1_ready         ( DownstreamStackBusLane[1][31].pe__std__lane_strm1_ready              ),      
        .std__pe1__lane31_strm1_cntl          ( DownstreamStackBusLane[1][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe1__lane31_strm1_data          ( DownstreamStackBusLane[1][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe1__lane31_strm1_data_valid    ( DownstreamStackBusLane[1][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane0_strm0_ready         ( DownstreamStackBusLane[2][0].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane0_strm0_cntl          ( DownstreamStackBusLane[2][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane0_strm0_data          ( DownstreamStackBusLane[2][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane0_strm0_data_valid    ( DownstreamStackBusLane[2][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane0_strm1_ready         ( DownstreamStackBusLane[2][0].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane0_strm1_cntl          ( DownstreamStackBusLane[2][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane0_strm1_data          ( DownstreamStackBusLane[2][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane0_strm1_data_valid    ( DownstreamStackBusLane[2][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane1_strm0_ready         ( DownstreamStackBusLane[2][1].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane1_strm0_cntl          ( DownstreamStackBusLane[2][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane1_strm0_data          ( DownstreamStackBusLane[2][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane1_strm0_data_valid    ( DownstreamStackBusLane[2][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane1_strm1_ready         ( DownstreamStackBusLane[2][1].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane1_strm1_cntl          ( DownstreamStackBusLane[2][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane1_strm1_data          ( DownstreamStackBusLane[2][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane1_strm1_data_valid    ( DownstreamStackBusLane[2][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane2_strm0_ready         ( DownstreamStackBusLane[2][2].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane2_strm0_cntl          ( DownstreamStackBusLane[2][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane2_strm0_data          ( DownstreamStackBusLane[2][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane2_strm0_data_valid    ( DownstreamStackBusLane[2][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane2_strm1_ready         ( DownstreamStackBusLane[2][2].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane2_strm1_cntl          ( DownstreamStackBusLane[2][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane2_strm1_data          ( DownstreamStackBusLane[2][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane2_strm1_data_valid    ( DownstreamStackBusLane[2][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane3_strm0_ready         ( DownstreamStackBusLane[2][3].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane3_strm0_cntl          ( DownstreamStackBusLane[2][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane3_strm0_data          ( DownstreamStackBusLane[2][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane3_strm0_data_valid    ( DownstreamStackBusLane[2][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane3_strm1_ready         ( DownstreamStackBusLane[2][3].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane3_strm1_cntl          ( DownstreamStackBusLane[2][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane3_strm1_data          ( DownstreamStackBusLane[2][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane3_strm1_data_valid    ( DownstreamStackBusLane[2][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane4_strm0_ready         ( DownstreamStackBusLane[2][4].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane4_strm0_cntl          ( DownstreamStackBusLane[2][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane4_strm0_data          ( DownstreamStackBusLane[2][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane4_strm0_data_valid    ( DownstreamStackBusLane[2][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane4_strm1_ready         ( DownstreamStackBusLane[2][4].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane4_strm1_cntl          ( DownstreamStackBusLane[2][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane4_strm1_data          ( DownstreamStackBusLane[2][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane4_strm1_data_valid    ( DownstreamStackBusLane[2][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane5_strm0_ready         ( DownstreamStackBusLane[2][5].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane5_strm0_cntl          ( DownstreamStackBusLane[2][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane5_strm0_data          ( DownstreamStackBusLane[2][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane5_strm0_data_valid    ( DownstreamStackBusLane[2][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane5_strm1_ready         ( DownstreamStackBusLane[2][5].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane5_strm1_cntl          ( DownstreamStackBusLane[2][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane5_strm1_data          ( DownstreamStackBusLane[2][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane5_strm1_data_valid    ( DownstreamStackBusLane[2][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane6_strm0_ready         ( DownstreamStackBusLane[2][6].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane6_strm0_cntl          ( DownstreamStackBusLane[2][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane6_strm0_data          ( DownstreamStackBusLane[2][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane6_strm0_data_valid    ( DownstreamStackBusLane[2][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane6_strm1_ready         ( DownstreamStackBusLane[2][6].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane6_strm1_cntl          ( DownstreamStackBusLane[2][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane6_strm1_data          ( DownstreamStackBusLane[2][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane6_strm1_data_valid    ( DownstreamStackBusLane[2][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane7_strm0_ready         ( DownstreamStackBusLane[2][7].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane7_strm0_cntl          ( DownstreamStackBusLane[2][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane7_strm0_data          ( DownstreamStackBusLane[2][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane7_strm0_data_valid    ( DownstreamStackBusLane[2][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane7_strm1_ready         ( DownstreamStackBusLane[2][7].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane7_strm1_cntl          ( DownstreamStackBusLane[2][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane7_strm1_data          ( DownstreamStackBusLane[2][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane7_strm1_data_valid    ( DownstreamStackBusLane[2][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane8_strm0_ready         ( DownstreamStackBusLane[2][8].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane8_strm0_cntl          ( DownstreamStackBusLane[2][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane8_strm0_data          ( DownstreamStackBusLane[2][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane8_strm0_data_valid    ( DownstreamStackBusLane[2][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane8_strm1_ready         ( DownstreamStackBusLane[2][8].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane8_strm1_cntl          ( DownstreamStackBusLane[2][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane8_strm1_data          ( DownstreamStackBusLane[2][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane8_strm1_data_valid    ( DownstreamStackBusLane[2][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane9_strm0_ready         ( DownstreamStackBusLane[2][9].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane9_strm0_cntl          ( DownstreamStackBusLane[2][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane9_strm0_data          ( DownstreamStackBusLane[2][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane9_strm0_data_valid    ( DownstreamStackBusLane[2][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane9_strm1_ready         ( DownstreamStackBusLane[2][9].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane9_strm1_cntl          ( DownstreamStackBusLane[2][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane9_strm1_data          ( DownstreamStackBusLane[2][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane9_strm1_data_valid    ( DownstreamStackBusLane[2][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane10_strm0_ready         ( DownstreamStackBusLane[2][10].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane10_strm0_cntl          ( DownstreamStackBusLane[2][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane10_strm0_data          ( DownstreamStackBusLane[2][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane10_strm0_data_valid    ( DownstreamStackBusLane[2][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane10_strm1_ready         ( DownstreamStackBusLane[2][10].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane10_strm1_cntl          ( DownstreamStackBusLane[2][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane10_strm1_data          ( DownstreamStackBusLane[2][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane10_strm1_data_valid    ( DownstreamStackBusLane[2][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane11_strm0_ready         ( DownstreamStackBusLane[2][11].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane11_strm0_cntl          ( DownstreamStackBusLane[2][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane11_strm0_data          ( DownstreamStackBusLane[2][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane11_strm0_data_valid    ( DownstreamStackBusLane[2][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane11_strm1_ready         ( DownstreamStackBusLane[2][11].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane11_strm1_cntl          ( DownstreamStackBusLane[2][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane11_strm1_data          ( DownstreamStackBusLane[2][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane11_strm1_data_valid    ( DownstreamStackBusLane[2][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane12_strm0_ready         ( DownstreamStackBusLane[2][12].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane12_strm0_cntl          ( DownstreamStackBusLane[2][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane12_strm0_data          ( DownstreamStackBusLane[2][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane12_strm0_data_valid    ( DownstreamStackBusLane[2][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane12_strm1_ready         ( DownstreamStackBusLane[2][12].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane12_strm1_cntl          ( DownstreamStackBusLane[2][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane12_strm1_data          ( DownstreamStackBusLane[2][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane12_strm1_data_valid    ( DownstreamStackBusLane[2][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane13_strm0_ready         ( DownstreamStackBusLane[2][13].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane13_strm0_cntl          ( DownstreamStackBusLane[2][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane13_strm0_data          ( DownstreamStackBusLane[2][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane13_strm0_data_valid    ( DownstreamStackBusLane[2][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane13_strm1_ready         ( DownstreamStackBusLane[2][13].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane13_strm1_cntl          ( DownstreamStackBusLane[2][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane13_strm1_data          ( DownstreamStackBusLane[2][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane13_strm1_data_valid    ( DownstreamStackBusLane[2][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane14_strm0_ready         ( DownstreamStackBusLane[2][14].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane14_strm0_cntl          ( DownstreamStackBusLane[2][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane14_strm0_data          ( DownstreamStackBusLane[2][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane14_strm0_data_valid    ( DownstreamStackBusLane[2][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane14_strm1_ready         ( DownstreamStackBusLane[2][14].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane14_strm1_cntl          ( DownstreamStackBusLane[2][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane14_strm1_data          ( DownstreamStackBusLane[2][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane14_strm1_data_valid    ( DownstreamStackBusLane[2][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane15_strm0_ready         ( DownstreamStackBusLane[2][15].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane15_strm0_cntl          ( DownstreamStackBusLane[2][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane15_strm0_data          ( DownstreamStackBusLane[2][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane15_strm0_data_valid    ( DownstreamStackBusLane[2][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane15_strm1_ready         ( DownstreamStackBusLane[2][15].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane15_strm1_cntl          ( DownstreamStackBusLane[2][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane15_strm1_data          ( DownstreamStackBusLane[2][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane15_strm1_data_valid    ( DownstreamStackBusLane[2][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane16_strm0_ready         ( DownstreamStackBusLane[2][16].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane16_strm0_cntl          ( DownstreamStackBusLane[2][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane16_strm0_data          ( DownstreamStackBusLane[2][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane16_strm0_data_valid    ( DownstreamStackBusLane[2][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane16_strm1_ready         ( DownstreamStackBusLane[2][16].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane16_strm1_cntl          ( DownstreamStackBusLane[2][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane16_strm1_data          ( DownstreamStackBusLane[2][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane16_strm1_data_valid    ( DownstreamStackBusLane[2][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane17_strm0_ready         ( DownstreamStackBusLane[2][17].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane17_strm0_cntl          ( DownstreamStackBusLane[2][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane17_strm0_data          ( DownstreamStackBusLane[2][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane17_strm0_data_valid    ( DownstreamStackBusLane[2][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane17_strm1_ready         ( DownstreamStackBusLane[2][17].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane17_strm1_cntl          ( DownstreamStackBusLane[2][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane17_strm1_data          ( DownstreamStackBusLane[2][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane17_strm1_data_valid    ( DownstreamStackBusLane[2][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane18_strm0_ready         ( DownstreamStackBusLane[2][18].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane18_strm0_cntl          ( DownstreamStackBusLane[2][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane18_strm0_data          ( DownstreamStackBusLane[2][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane18_strm0_data_valid    ( DownstreamStackBusLane[2][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane18_strm1_ready         ( DownstreamStackBusLane[2][18].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane18_strm1_cntl          ( DownstreamStackBusLane[2][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane18_strm1_data          ( DownstreamStackBusLane[2][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane18_strm1_data_valid    ( DownstreamStackBusLane[2][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane19_strm0_ready         ( DownstreamStackBusLane[2][19].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane19_strm0_cntl          ( DownstreamStackBusLane[2][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane19_strm0_data          ( DownstreamStackBusLane[2][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane19_strm0_data_valid    ( DownstreamStackBusLane[2][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane19_strm1_ready         ( DownstreamStackBusLane[2][19].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane19_strm1_cntl          ( DownstreamStackBusLane[2][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane19_strm1_data          ( DownstreamStackBusLane[2][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane19_strm1_data_valid    ( DownstreamStackBusLane[2][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane20_strm0_ready         ( DownstreamStackBusLane[2][20].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane20_strm0_cntl          ( DownstreamStackBusLane[2][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane20_strm0_data          ( DownstreamStackBusLane[2][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane20_strm0_data_valid    ( DownstreamStackBusLane[2][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane20_strm1_ready         ( DownstreamStackBusLane[2][20].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane20_strm1_cntl          ( DownstreamStackBusLane[2][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane20_strm1_data          ( DownstreamStackBusLane[2][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane20_strm1_data_valid    ( DownstreamStackBusLane[2][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane21_strm0_ready         ( DownstreamStackBusLane[2][21].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane21_strm0_cntl          ( DownstreamStackBusLane[2][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane21_strm0_data          ( DownstreamStackBusLane[2][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane21_strm0_data_valid    ( DownstreamStackBusLane[2][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane21_strm1_ready         ( DownstreamStackBusLane[2][21].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane21_strm1_cntl          ( DownstreamStackBusLane[2][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane21_strm1_data          ( DownstreamStackBusLane[2][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane21_strm1_data_valid    ( DownstreamStackBusLane[2][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane22_strm0_ready         ( DownstreamStackBusLane[2][22].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane22_strm0_cntl          ( DownstreamStackBusLane[2][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane22_strm0_data          ( DownstreamStackBusLane[2][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane22_strm0_data_valid    ( DownstreamStackBusLane[2][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane22_strm1_ready         ( DownstreamStackBusLane[2][22].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane22_strm1_cntl          ( DownstreamStackBusLane[2][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane22_strm1_data          ( DownstreamStackBusLane[2][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane22_strm1_data_valid    ( DownstreamStackBusLane[2][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane23_strm0_ready         ( DownstreamStackBusLane[2][23].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane23_strm0_cntl          ( DownstreamStackBusLane[2][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane23_strm0_data          ( DownstreamStackBusLane[2][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane23_strm0_data_valid    ( DownstreamStackBusLane[2][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane23_strm1_ready         ( DownstreamStackBusLane[2][23].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane23_strm1_cntl          ( DownstreamStackBusLane[2][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane23_strm1_data          ( DownstreamStackBusLane[2][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane23_strm1_data_valid    ( DownstreamStackBusLane[2][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane24_strm0_ready         ( DownstreamStackBusLane[2][24].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane24_strm0_cntl          ( DownstreamStackBusLane[2][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane24_strm0_data          ( DownstreamStackBusLane[2][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane24_strm0_data_valid    ( DownstreamStackBusLane[2][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane24_strm1_ready         ( DownstreamStackBusLane[2][24].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane24_strm1_cntl          ( DownstreamStackBusLane[2][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane24_strm1_data          ( DownstreamStackBusLane[2][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane24_strm1_data_valid    ( DownstreamStackBusLane[2][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane25_strm0_ready         ( DownstreamStackBusLane[2][25].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane25_strm0_cntl          ( DownstreamStackBusLane[2][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane25_strm0_data          ( DownstreamStackBusLane[2][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane25_strm0_data_valid    ( DownstreamStackBusLane[2][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane25_strm1_ready         ( DownstreamStackBusLane[2][25].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane25_strm1_cntl          ( DownstreamStackBusLane[2][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane25_strm1_data          ( DownstreamStackBusLane[2][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane25_strm1_data_valid    ( DownstreamStackBusLane[2][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane26_strm0_ready         ( DownstreamStackBusLane[2][26].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane26_strm0_cntl          ( DownstreamStackBusLane[2][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane26_strm0_data          ( DownstreamStackBusLane[2][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane26_strm0_data_valid    ( DownstreamStackBusLane[2][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane26_strm1_ready         ( DownstreamStackBusLane[2][26].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane26_strm1_cntl          ( DownstreamStackBusLane[2][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane26_strm1_data          ( DownstreamStackBusLane[2][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane26_strm1_data_valid    ( DownstreamStackBusLane[2][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane27_strm0_ready         ( DownstreamStackBusLane[2][27].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane27_strm0_cntl          ( DownstreamStackBusLane[2][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane27_strm0_data          ( DownstreamStackBusLane[2][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane27_strm0_data_valid    ( DownstreamStackBusLane[2][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane27_strm1_ready         ( DownstreamStackBusLane[2][27].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane27_strm1_cntl          ( DownstreamStackBusLane[2][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane27_strm1_data          ( DownstreamStackBusLane[2][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane27_strm1_data_valid    ( DownstreamStackBusLane[2][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane28_strm0_ready         ( DownstreamStackBusLane[2][28].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane28_strm0_cntl          ( DownstreamStackBusLane[2][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane28_strm0_data          ( DownstreamStackBusLane[2][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane28_strm0_data_valid    ( DownstreamStackBusLane[2][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane28_strm1_ready         ( DownstreamStackBusLane[2][28].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane28_strm1_cntl          ( DownstreamStackBusLane[2][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane28_strm1_data          ( DownstreamStackBusLane[2][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane28_strm1_data_valid    ( DownstreamStackBusLane[2][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane29_strm0_ready         ( DownstreamStackBusLane[2][29].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane29_strm0_cntl          ( DownstreamStackBusLane[2][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane29_strm0_data          ( DownstreamStackBusLane[2][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane29_strm0_data_valid    ( DownstreamStackBusLane[2][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane29_strm1_ready         ( DownstreamStackBusLane[2][29].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane29_strm1_cntl          ( DownstreamStackBusLane[2][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane29_strm1_data          ( DownstreamStackBusLane[2][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane29_strm1_data_valid    ( DownstreamStackBusLane[2][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane30_strm0_ready         ( DownstreamStackBusLane[2][30].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane30_strm0_cntl          ( DownstreamStackBusLane[2][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane30_strm0_data          ( DownstreamStackBusLane[2][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane30_strm0_data_valid    ( DownstreamStackBusLane[2][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane30_strm1_ready         ( DownstreamStackBusLane[2][30].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane30_strm1_cntl          ( DownstreamStackBusLane[2][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane30_strm1_data          ( DownstreamStackBusLane[2][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane30_strm1_data_valid    ( DownstreamStackBusLane[2][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 2, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane31_strm0_ready         ( DownstreamStackBusLane[2][31].pe__std__lane_strm0_ready              ),      
        .std__pe2__lane31_strm0_cntl          ( DownstreamStackBusLane[2][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe2__lane31_strm0_data          ( DownstreamStackBusLane[2][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe2__lane31_strm0_data_valid    ( DownstreamStackBusLane[2][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__std__lane31_strm1_ready         ( DownstreamStackBusLane[2][31].pe__std__lane_strm1_ready              ),      
        .std__pe2__lane31_strm1_cntl          ( DownstreamStackBusLane[2][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe2__lane31_strm1_data          ( DownstreamStackBusLane[2][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe2__lane31_strm1_data_valid    ( DownstreamStackBusLane[2][31].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane0_strm0_ready         ( DownstreamStackBusLane[3][0].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane0_strm0_cntl          ( DownstreamStackBusLane[3][0].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane0_strm0_data          ( DownstreamStackBusLane[3][0].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane0_strm0_data_valid    ( DownstreamStackBusLane[3][0].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane0_strm1_ready         ( DownstreamStackBusLane[3][0].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane0_strm1_cntl          ( DownstreamStackBusLane[3][0].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane0_strm1_data          ( DownstreamStackBusLane[3][0].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane0_strm1_data_valid    ( DownstreamStackBusLane[3][0].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane1_strm0_ready         ( DownstreamStackBusLane[3][1].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane1_strm0_cntl          ( DownstreamStackBusLane[3][1].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane1_strm0_data          ( DownstreamStackBusLane[3][1].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane1_strm0_data_valid    ( DownstreamStackBusLane[3][1].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane1_strm1_ready         ( DownstreamStackBusLane[3][1].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane1_strm1_cntl          ( DownstreamStackBusLane[3][1].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane1_strm1_data          ( DownstreamStackBusLane[3][1].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane1_strm1_data_valid    ( DownstreamStackBusLane[3][1].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane2_strm0_ready         ( DownstreamStackBusLane[3][2].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane2_strm0_cntl          ( DownstreamStackBusLane[3][2].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane2_strm0_data          ( DownstreamStackBusLane[3][2].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane2_strm0_data_valid    ( DownstreamStackBusLane[3][2].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane2_strm1_ready         ( DownstreamStackBusLane[3][2].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane2_strm1_cntl          ( DownstreamStackBusLane[3][2].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane2_strm1_data          ( DownstreamStackBusLane[3][2].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane2_strm1_data_valid    ( DownstreamStackBusLane[3][2].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane3_strm0_ready         ( DownstreamStackBusLane[3][3].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane3_strm0_cntl          ( DownstreamStackBusLane[3][3].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane3_strm0_data          ( DownstreamStackBusLane[3][3].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane3_strm0_data_valid    ( DownstreamStackBusLane[3][3].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane3_strm1_ready         ( DownstreamStackBusLane[3][3].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane3_strm1_cntl          ( DownstreamStackBusLane[3][3].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane3_strm1_data          ( DownstreamStackBusLane[3][3].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane3_strm1_data_valid    ( DownstreamStackBusLane[3][3].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane4_strm0_ready         ( DownstreamStackBusLane[3][4].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane4_strm0_cntl          ( DownstreamStackBusLane[3][4].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane4_strm0_data          ( DownstreamStackBusLane[3][4].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane4_strm0_data_valid    ( DownstreamStackBusLane[3][4].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane4_strm1_ready         ( DownstreamStackBusLane[3][4].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane4_strm1_cntl          ( DownstreamStackBusLane[3][4].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane4_strm1_data          ( DownstreamStackBusLane[3][4].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane4_strm1_data_valid    ( DownstreamStackBusLane[3][4].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane5_strm0_ready         ( DownstreamStackBusLane[3][5].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane5_strm0_cntl          ( DownstreamStackBusLane[3][5].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane5_strm0_data          ( DownstreamStackBusLane[3][5].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane5_strm0_data_valid    ( DownstreamStackBusLane[3][5].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane5_strm1_ready         ( DownstreamStackBusLane[3][5].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane5_strm1_cntl          ( DownstreamStackBusLane[3][5].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane5_strm1_data          ( DownstreamStackBusLane[3][5].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane5_strm1_data_valid    ( DownstreamStackBusLane[3][5].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane6_strm0_ready         ( DownstreamStackBusLane[3][6].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane6_strm0_cntl          ( DownstreamStackBusLane[3][6].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane6_strm0_data          ( DownstreamStackBusLane[3][6].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane6_strm0_data_valid    ( DownstreamStackBusLane[3][6].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane6_strm1_ready         ( DownstreamStackBusLane[3][6].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane6_strm1_cntl          ( DownstreamStackBusLane[3][6].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane6_strm1_data          ( DownstreamStackBusLane[3][6].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane6_strm1_data_valid    ( DownstreamStackBusLane[3][6].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane7_strm0_ready         ( DownstreamStackBusLane[3][7].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane7_strm0_cntl          ( DownstreamStackBusLane[3][7].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane7_strm0_data          ( DownstreamStackBusLane[3][7].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane7_strm0_data_valid    ( DownstreamStackBusLane[3][7].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane7_strm1_ready         ( DownstreamStackBusLane[3][7].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane7_strm1_cntl          ( DownstreamStackBusLane[3][7].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane7_strm1_data          ( DownstreamStackBusLane[3][7].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane7_strm1_data_valid    ( DownstreamStackBusLane[3][7].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane8_strm0_ready         ( DownstreamStackBusLane[3][8].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane8_strm0_cntl          ( DownstreamStackBusLane[3][8].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane8_strm0_data          ( DownstreamStackBusLane[3][8].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane8_strm0_data_valid    ( DownstreamStackBusLane[3][8].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane8_strm1_ready         ( DownstreamStackBusLane[3][8].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane8_strm1_cntl          ( DownstreamStackBusLane[3][8].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane8_strm1_data          ( DownstreamStackBusLane[3][8].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane8_strm1_data_valid    ( DownstreamStackBusLane[3][8].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane9_strm0_ready         ( DownstreamStackBusLane[3][9].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane9_strm0_cntl          ( DownstreamStackBusLane[3][9].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane9_strm0_data          ( DownstreamStackBusLane[3][9].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane9_strm0_data_valid    ( DownstreamStackBusLane[3][9].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane9_strm1_ready         ( DownstreamStackBusLane[3][9].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane9_strm1_cntl          ( DownstreamStackBusLane[3][9].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane9_strm1_data          ( DownstreamStackBusLane[3][9].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane9_strm1_data_valid    ( DownstreamStackBusLane[3][9].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane10_strm0_ready         ( DownstreamStackBusLane[3][10].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane10_strm0_cntl          ( DownstreamStackBusLane[3][10].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane10_strm0_data          ( DownstreamStackBusLane[3][10].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane10_strm0_data_valid    ( DownstreamStackBusLane[3][10].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane10_strm1_ready         ( DownstreamStackBusLane[3][10].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane10_strm1_cntl          ( DownstreamStackBusLane[3][10].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane10_strm1_data          ( DownstreamStackBusLane[3][10].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane10_strm1_data_valid    ( DownstreamStackBusLane[3][10].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane11_strm0_ready         ( DownstreamStackBusLane[3][11].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane11_strm0_cntl          ( DownstreamStackBusLane[3][11].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane11_strm0_data          ( DownstreamStackBusLane[3][11].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane11_strm0_data_valid    ( DownstreamStackBusLane[3][11].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane11_strm1_ready         ( DownstreamStackBusLane[3][11].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane11_strm1_cntl          ( DownstreamStackBusLane[3][11].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane11_strm1_data          ( DownstreamStackBusLane[3][11].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane11_strm1_data_valid    ( DownstreamStackBusLane[3][11].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane12_strm0_ready         ( DownstreamStackBusLane[3][12].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane12_strm0_cntl          ( DownstreamStackBusLane[3][12].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane12_strm0_data          ( DownstreamStackBusLane[3][12].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane12_strm0_data_valid    ( DownstreamStackBusLane[3][12].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane12_strm1_ready         ( DownstreamStackBusLane[3][12].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane12_strm1_cntl          ( DownstreamStackBusLane[3][12].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane12_strm1_data          ( DownstreamStackBusLane[3][12].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane12_strm1_data_valid    ( DownstreamStackBusLane[3][12].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane13_strm0_ready         ( DownstreamStackBusLane[3][13].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane13_strm0_cntl          ( DownstreamStackBusLane[3][13].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane13_strm0_data          ( DownstreamStackBusLane[3][13].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane13_strm0_data_valid    ( DownstreamStackBusLane[3][13].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane13_strm1_ready         ( DownstreamStackBusLane[3][13].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane13_strm1_cntl          ( DownstreamStackBusLane[3][13].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane13_strm1_data          ( DownstreamStackBusLane[3][13].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane13_strm1_data_valid    ( DownstreamStackBusLane[3][13].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane14_strm0_ready         ( DownstreamStackBusLane[3][14].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane14_strm0_cntl          ( DownstreamStackBusLane[3][14].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane14_strm0_data          ( DownstreamStackBusLane[3][14].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane14_strm0_data_valid    ( DownstreamStackBusLane[3][14].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane14_strm1_ready         ( DownstreamStackBusLane[3][14].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane14_strm1_cntl          ( DownstreamStackBusLane[3][14].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane14_strm1_data          ( DownstreamStackBusLane[3][14].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane14_strm1_data_valid    ( DownstreamStackBusLane[3][14].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane15_strm0_ready         ( DownstreamStackBusLane[3][15].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane15_strm0_cntl          ( DownstreamStackBusLane[3][15].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane15_strm0_data          ( DownstreamStackBusLane[3][15].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane15_strm0_data_valid    ( DownstreamStackBusLane[3][15].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane15_strm1_ready         ( DownstreamStackBusLane[3][15].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane15_strm1_cntl          ( DownstreamStackBusLane[3][15].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane15_strm1_data          ( DownstreamStackBusLane[3][15].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane15_strm1_data_valid    ( DownstreamStackBusLane[3][15].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane16_strm0_ready         ( DownstreamStackBusLane[3][16].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane16_strm0_cntl          ( DownstreamStackBusLane[3][16].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane16_strm0_data          ( DownstreamStackBusLane[3][16].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane16_strm0_data_valid    ( DownstreamStackBusLane[3][16].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane16_strm1_ready         ( DownstreamStackBusLane[3][16].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane16_strm1_cntl          ( DownstreamStackBusLane[3][16].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane16_strm1_data          ( DownstreamStackBusLane[3][16].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane16_strm1_data_valid    ( DownstreamStackBusLane[3][16].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane17_strm0_ready         ( DownstreamStackBusLane[3][17].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane17_strm0_cntl          ( DownstreamStackBusLane[3][17].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane17_strm0_data          ( DownstreamStackBusLane[3][17].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane17_strm0_data_valid    ( DownstreamStackBusLane[3][17].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane17_strm1_ready         ( DownstreamStackBusLane[3][17].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane17_strm1_cntl          ( DownstreamStackBusLane[3][17].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane17_strm1_data          ( DownstreamStackBusLane[3][17].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane17_strm1_data_valid    ( DownstreamStackBusLane[3][17].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane18_strm0_ready         ( DownstreamStackBusLane[3][18].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane18_strm0_cntl          ( DownstreamStackBusLane[3][18].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane18_strm0_data          ( DownstreamStackBusLane[3][18].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane18_strm0_data_valid    ( DownstreamStackBusLane[3][18].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane18_strm1_ready         ( DownstreamStackBusLane[3][18].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane18_strm1_cntl          ( DownstreamStackBusLane[3][18].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane18_strm1_data          ( DownstreamStackBusLane[3][18].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane18_strm1_data_valid    ( DownstreamStackBusLane[3][18].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane19_strm0_ready         ( DownstreamStackBusLane[3][19].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane19_strm0_cntl          ( DownstreamStackBusLane[3][19].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane19_strm0_data          ( DownstreamStackBusLane[3][19].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane19_strm0_data_valid    ( DownstreamStackBusLane[3][19].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane19_strm1_ready         ( DownstreamStackBusLane[3][19].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane19_strm1_cntl          ( DownstreamStackBusLane[3][19].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane19_strm1_data          ( DownstreamStackBusLane[3][19].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane19_strm1_data_valid    ( DownstreamStackBusLane[3][19].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane20_strm0_ready         ( DownstreamStackBusLane[3][20].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane20_strm0_cntl          ( DownstreamStackBusLane[3][20].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane20_strm0_data          ( DownstreamStackBusLane[3][20].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane20_strm0_data_valid    ( DownstreamStackBusLane[3][20].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane20_strm1_ready         ( DownstreamStackBusLane[3][20].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane20_strm1_cntl          ( DownstreamStackBusLane[3][20].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane20_strm1_data          ( DownstreamStackBusLane[3][20].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane20_strm1_data_valid    ( DownstreamStackBusLane[3][20].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane21_strm0_ready         ( DownstreamStackBusLane[3][21].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane21_strm0_cntl          ( DownstreamStackBusLane[3][21].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane21_strm0_data          ( DownstreamStackBusLane[3][21].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane21_strm0_data_valid    ( DownstreamStackBusLane[3][21].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane21_strm1_ready         ( DownstreamStackBusLane[3][21].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane21_strm1_cntl          ( DownstreamStackBusLane[3][21].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane21_strm1_data          ( DownstreamStackBusLane[3][21].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane21_strm1_data_valid    ( DownstreamStackBusLane[3][21].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane22_strm0_ready         ( DownstreamStackBusLane[3][22].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane22_strm0_cntl          ( DownstreamStackBusLane[3][22].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane22_strm0_data          ( DownstreamStackBusLane[3][22].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane22_strm0_data_valid    ( DownstreamStackBusLane[3][22].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane22_strm1_ready         ( DownstreamStackBusLane[3][22].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane22_strm1_cntl          ( DownstreamStackBusLane[3][22].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane22_strm1_data          ( DownstreamStackBusLane[3][22].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane22_strm1_data_valid    ( DownstreamStackBusLane[3][22].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane23_strm0_ready         ( DownstreamStackBusLane[3][23].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane23_strm0_cntl          ( DownstreamStackBusLane[3][23].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane23_strm0_data          ( DownstreamStackBusLane[3][23].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane23_strm0_data_valid    ( DownstreamStackBusLane[3][23].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane23_strm1_ready         ( DownstreamStackBusLane[3][23].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane23_strm1_cntl          ( DownstreamStackBusLane[3][23].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane23_strm1_data          ( DownstreamStackBusLane[3][23].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane23_strm1_data_valid    ( DownstreamStackBusLane[3][23].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane24_strm0_ready         ( DownstreamStackBusLane[3][24].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane24_strm0_cntl          ( DownstreamStackBusLane[3][24].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane24_strm0_data          ( DownstreamStackBusLane[3][24].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane24_strm0_data_valid    ( DownstreamStackBusLane[3][24].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane24_strm1_ready         ( DownstreamStackBusLane[3][24].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane24_strm1_cntl          ( DownstreamStackBusLane[3][24].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane24_strm1_data          ( DownstreamStackBusLane[3][24].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane24_strm1_data_valid    ( DownstreamStackBusLane[3][24].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane25_strm0_ready         ( DownstreamStackBusLane[3][25].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane25_strm0_cntl          ( DownstreamStackBusLane[3][25].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane25_strm0_data          ( DownstreamStackBusLane[3][25].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane25_strm0_data_valid    ( DownstreamStackBusLane[3][25].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane25_strm1_ready         ( DownstreamStackBusLane[3][25].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane25_strm1_cntl          ( DownstreamStackBusLane[3][25].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane25_strm1_data          ( DownstreamStackBusLane[3][25].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane25_strm1_data_valid    ( DownstreamStackBusLane[3][25].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane26_strm0_ready         ( DownstreamStackBusLane[3][26].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane26_strm0_cntl          ( DownstreamStackBusLane[3][26].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane26_strm0_data          ( DownstreamStackBusLane[3][26].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane26_strm0_data_valid    ( DownstreamStackBusLane[3][26].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane26_strm1_ready         ( DownstreamStackBusLane[3][26].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane26_strm1_cntl          ( DownstreamStackBusLane[3][26].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane26_strm1_data          ( DownstreamStackBusLane[3][26].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane26_strm1_data_valid    ( DownstreamStackBusLane[3][26].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane27_strm0_ready         ( DownstreamStackBusLane[3][27].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane27_strm0_cntl          ( DownstreamStackBusLane[3][27].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane27_strm0_data          ( DownstreamStackBusLane[3][27].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane27_strm0_data_valid    ( DownstreamStackBusLane[3][27].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane27_strm1_ready         ( DownstreamStackBusLane[3][27].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane27_strm1_cntl          ( DownstreamStackBusLane[3][27].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane27_strm1_data          ( DownstreamStackBusLane[3][27].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane27_strm1_data_valid    ( DownstreamStackBusLane[3][27].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane28_strm0_ready         ( DownstreamStackBusLane[3][28].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane28_strm0_cntl          ( DownstreamStackBusLane[3][28].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane28_strm0_data          ( DownstreamStackBusLane[3][28].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane28_strm0_data_valid    ( DownstreamStackBusLane[3][28].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane28_strm1_ready         ( DownstreamStackBusLane[3][28].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane28_strm1_cntl          ( DownstreamStackBusLane[3][28].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane28_strm1_data          ( DownstreamStackBusLane[3][28].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane28_strm1_data_valid    ( DownstreamStackBusLane[3][28].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane29_strm0_ready         ( DownstreamStackBusLane[3][29].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane29_strm0_cntl          ( DownstreamStackBusLane[3][29].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane29_strm0_data          ( DownstreamStackBusLane[3][29].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane29_strm0_data_valid    ( DownstreamStackBusLane[3][29].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane29_strm1_ready         ( DownstreamStackBusLane[3][29].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane29_strm1_cntl          ( DownstreamStackBusLane[3][29].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane29_strm1_data          ( DownstreamStackBusLane[3][29].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane29_strm1_data_valid    ( DownstreamStackBusLane[3][29].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane30_strm0_ready         ( DownstreamStackBusLane[3][30].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane30_strm0_cntl          ( DownstreamStackBusLane[3][30].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane30_strm0_data          ( DownstreamStackBusLane[3][30].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane30_strm0_data_valid    ( DownstreamStackBusLane[3][30].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane30_strm1_ready         ( DownstreamStackBusLane[3][30].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane30_strm1_cntl          ( DownstreamStackBusLane[3][30].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane30_strm1_data          ( DownstreamStackBusLane[3][30].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane30_strm1_data_valid    ( DownstreamStackBusLane[3][30].cb_test.std__pe__lane_strm1_data_valid ),      
        
        // PE 3, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane31_strm0_ready         ( DownstreamStackBusLane[3][31].pe__std__lane_strm0_ready              ),      
        .std__pe3__lane31_strm0_cntl          ( DownstreamStackBusLane[3][31].cb_test.std__pe__lane_strm0_cntl       ),      
        .std__pe3__lane31_strm0_data          ( DownstreamStackBusLane[3][31].cb_test.std__pe__lane_strm0_data       ),      
        .std__pe3__lane31_strm0_data_valid    ( DownstreamStackBusLane[3][31].cb_test.std__pe__lane_strm0_data_valid ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__std__lane31_strm1_ready         ( DownstreamStackBusLane[3][31].pe__std__lane_strm1_ready              ),      
        .std__pe3__lane31_strm1_cntl          ( DownstreamStackBusLane[3][31].cb_test.std__pe__lane_strm1_cntl       ),      
        .std__pe3__lane31_strm1_data          ( DownstreamStackBusLane[3][31].cb_test.std__pe__lane_strm1_data       ),      
        .std__pe3__lane31_strm1_data_valid    ( DownstreamStackBusLane[3][31].cb_test.std__pe__lane_strm1_data_valid ),      
        