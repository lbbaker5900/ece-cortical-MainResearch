`ifndef _manager_vh
`define _manager_vh

/*****************************************************************

    File name   : manager.vh
    Author      : Lee Baker
    Affiliation : North Carolina State University, Raleigh, NC
    Date        : Mar 2017
    email       : lbbaker@ncsu.edu

*****************************************************************/

//------------------------------------------------
// System
//------------------------------------------------
`define MGR_MGR_ID_WIDTH             (`CLOG2(`MGR_ARRAY_NUM_OF_MGR))
`define MGR_MGR_ID_MSB               (`MGR_MGR_ID_WIDTH-1)
`define MGR_MGR_ID_LSB               0
`define MGR_MGR_ID_SIZE              (`MGR_MGR_ID_MSB - `MGR_MGR_ID_LSB +1)
`define MGR_MGR_ID_RANGE              `MGR_MGR_ID_MSB : `MGR_MGR_ID_LSB

`define MGR_MGR_ID_BITMASK_WIDTH             `MGR_ARRAY_NUM_OF_MGR
`define MGR_MGR_ID_BITMASK_MSB               (`MGR_MGR_ID_BITMASK_WIDTH-1)
`define MGR_MGR_ID_BITMASK_LSB               0
`define MGR_MGR_ID_BITMASK_SIZE              (`MGR_MGR_ID_BITMASK_MSB - `MGR_MGR_ID_BITMASK_LSB +1)
`define MGR_MGR_ID_BITMASK_RANGE              `MGR_MGR_ID_BITMASK_MSB : `MGR_MGR_ID_BITMASK_LSB
//------------------------------------------------
// Stack Bus stream
//------------------------------------------------

// we will carry a tag to track result (to possibly support multiple operations before first result is returned)
`define MGR_STD_OOB_TAG_WIDTH          `PE_STD_OOB_TAG_WIDTH
`define MGR_STD_OOB_TAG_MSB            `MGR_STD_OOB_TAG_WIDTH-1
`define MGR_STD_OOB_TAG_LSB            0
`define MGR_STD_OOB_TAG_RANGE          `MGR_STD_OOB_TAG_MSB : `MGR_STD_OOB_TAG_LSB

`define MGR_STD_LANE_DATA_WIDTH          `STACK_DOWN_INTF_STRM_DATA_WIDTH 
`define MGR_STD_LANE_DATA_MSB            `MGR_STD_LANE_DATA_WIDTH-1
`define MGR_STD_LANE_DATA_LSB            0
`define MGR_STD_LANE_DATA_RANGE          `MGR_STD_LANE_DATA_MSB : `MGR_STD_LANE_DATA_LSB

`define MGR_STU_DATA_WIDTH          `STACK_UP_INTF_DATA_WIDTH 
`define MGR_STU_DATA_MSB            `MGR_STU_DATA_WIDTH-1
`define MGR_STU_DATA_LSB            0
`define MGR_STU_DATA_RANGE          `MGR_STU_DATA_MSB : `MGR_STU_DATA_LSB



//------------------------------------------------
// MGR Stack bus streams
//------------------------------------------------

`define MGR_NUM_OF_STREAMS               `PE_NUM_OF_STREAMS 
`define MGR_NUM_OF_STREAMS_MSB           (`MGR_NUM_OF_STREAMS -1)
`define MGR_NUM_OF_STREAMS_LSB            0
`define MGR_NUM_OF_STREAMS_SIZE           (`MGR_NUM_OF_STREAMS_MSB - `MGR_NUM_OF_STREAMS_LSB +1)
`define MGR_NUM_OF_STREAMS_RANGE           `MGR_NUM_OF_STREAMS_MSB : `MGR_NUM_OF_STREAMS_LSB

//------------------------------------------------
// MGR Execution Lane 
//------------------------------------------------

`define MGR_NUM_OF_EXEC_LANES               `PE_NUM_OF_EXEC_LANES
`define MGR_NUM_OF_EXEC_LANES_MSB           (`MGR_NUM_OF_EXEC_LANES -1)
`define MGR_NUM_OF_EXEC_LANES_LSB            0
`define MGR_NUM_OF_EXEC_LANES_SIZE           (`MGR_NUM_OF_EXEC_LANES_MSB - `MGR_NUM_OF_EXEC_LANES_LSB +1)
`define MGR_NUM_OF_EXEC_LANES_RANGE           `MGR_NUM_OF_EXEC_LANES_MSB : `MGR_NUM_OF_EXEC_LANES_LSB

`define MGR_EXEC_LANE_WIDTH               `PE_EXEC_LANE_WIDTH
`define MGR_EXEC_LANE_WIDTH_MSB           `MGR_EXEC_LANE_WIDTH-1
`define MGR_EXEC_LANE_WIDTH_LSB            0
`define MGR_EXEC_LANE_WIDTH_SIZE           (`MGR_EXEC_LANE_WIDTH_MSB - `MGR_EXEC_LANE_WIDTH_LSB +1)
`define MGR_EXEC_LANE_WIDTH_RANGE           `MGR_EXEC_LANE_WIDTH_MSB : `MGR_EXEC_LANE_WIDTH_LSB

`define MGR_EXEC_LANE_ID_WIDTH            `PE_EXEC_LANE_ID_WIDTH   
`define MGR_EXEC_LANE_ID_MSB              `PE_EXEC_LANE_ID_MSB     
`define MGR_EXEC_LANE_ID_LSB              `PE_EXEC_LANE_ID_LSB     
`define MGR_EXEC_LANE_ID_RANGE            `PE_EXEC_LANE_ID_RANGE   

//--------------------------------------------------------
// In cases where we set number of active lanes, Number of active lanes is 1..32, so need 6 bits
  
`define MGR_NUM_LANES_WIDTH               (`CLOG2(`PE_NUM_OF_EXEC_LANES))+1
`define MGR_NUM_LANES_MSB           `MGR_NUM_LANES_WIDTH-1
`define MGR_NUM_LANES_LSB            0
`define MGR_NUM_LANES_SIZE           (`MGR_NUM_LANES_MSB - `MGR_NUM_LANES_LSB +1)
`define MGR_NUM_LANES_RANGE           `MGR_NUM_LANES_MSB : `MGR_NUM_LANES_LSB
//---------------------------------------------------------------------------------------------------------------------
// Memory

//---------------------------------------------------------------------------------------------------------------------
// WU Memory

// FIXME
`define MGR_WU_MEMORY_DEPTH                      4096
`define MGR_WU_ADDRESS_WIDTH                       (`CLOG2(`MGR_WU_MEMORY_DEPTH))
`define MGR_WU_ADDRESS_MSB                         `MGR_WU_ADDRESS_WIDTH-1
`define MGR_WU_ADDRESS_LSB                         0
`define MGR_WU_ADDRESS_SIZE                        (`MGR_WU_ADDRESS_MSB - `MGR_WU_ADDRESS_LSB +1)
`define MGR_WU_ADDRESS_RANGE                        `MGR_WU_ADDRESS_MSB : `MGR_WU_ADDRESS_LSB



//---------------------------------------------------------------------------------------------------------------------
// WU Instruction

`define MGR_WU_OPT_PER_INST                       3
`define MGR_WU_OPT_PER_INST_WIDTH                 `MGR_WU_OPT_PER_INST   
`define MGR_WU_OPT_PER_INST_MSB                   `MGR_WU_OPT_PER_INST_WIDTH-1
`define MGR_WU_OPT_PER_INST_LSB                   0
`define MGR_WU_OPT_PER_INST_SIZE                  (`MGR_WU_OPT_PER_INST_MSB - `MGR_WU_OPT_PER_INST_LSB +1)
`define MGR_WU_OPT_PER_INST_RANGE                  `MGR_WU_OPT_PER_INST_MSB : `MGR_WU_OPT_PER_INST_LSB


`define MGR_WU_OPT_TYPE_WIDTH                 8
`define MGR_WU_OPT_TYPE_MSB                   `MGR_WU_OPT_TYPE_WIDTH-1
`define MGR_WU_OPT_TYPE_LSB                   0
`define MGR_WU_OPT_TYPE_SIZE                  (`MGR_WU_OPT_TYPE_MSB - `MGR_WU_OPT_TYPE_LSB +1)
`define MGR_WU_OPT_TYPE_RANGE                  `MGR_WU_OPT_TYPE_MSB : `MGR_WU_OPT_TYPE_LSB


`define MGR_WU_OPT_VALUE_WIDTH                 8
`define MGR_WU_OPT_VALUE_MSB                   `MGR_WU_OPT_VALUE_WIDTH-1
`define MGR_WU_OPT_VALUE_LSB                   0
`define MGR_WU_OPT_VALUE_SIZE                  (`MGR_WU_OPT_VALUE_MSB - `MGR_WU_OPT_VALUE_LSB +1)
`define MGR_WU_OPT_VALUE_RANGE                  `MGR_WU_OPT_VALUE_MSB : `MGR_WU_OPT_VALUE_LSB


`define MGR_WU_EXTD_OPT_VALUE_WIDTH                 `MGR_WU_OPT_VALUE_WIDTH  *3
`define MGR_WU_EXTD_OPT_VALUE_MSB                   `MGR_WU_EXTD_OPT_VALUE_WIDTH-1
`define MGR_WU_EXTD_OPT_VALUE_LSB                   0
`define MGR_WU_EXTD_OPT_VALUE_SIZE                  (`MGR_WU_EXTD_OPT_VALUE_MSB - `MGR_WU_EXTD_OPT_VALUE_LSB +1)
`define MGR_WU_EXTD_OPT_VALUE_RANGE                  `MGR_WU_EXTD_OPT_VALUE_MSB : `MGR_WU_EXTD_OPT_VALUE_LSB

`define MGR_WU_TUPLE_WIDTH                 'MGR_WU_OPT_TYPE_WIDTH+`MGR_WU_OPT_VALUE_WIDTH
`define MGR_WU_TUPLE_MSB                   `MGR_WU_TUPLE_WIDTH-1
`define MGR_WU_TUPLE_LSB                   0
`define MGR_WU_TUPLE_SIZE                  (`MGR_WU_TUPLE_MSB - `MGR_WU_TUPLE_LSB +1)
`define MGR_WU_TUPLE_RANGE                  `MGR_WU_TUPLE_MSB : `MGR_WU_TUPLE_LSB

`define MGR_WU_EXTD_TUPLE_WIDTH            'MGR_WU_OPT_TYPE_WIDTH+`MGR_WU_EXTD_OPT_VALUE_WIDTH
`define MGR_WU_EXTD_TUPLE_MSB              `MGR_WU_EXTD_TUPLE_WIDTH-1
`define MGR_WU_EXTD_TUPLE_LSB              0
`define MGR_WU_EXTD_TUPLE_SIZE             (`MGR_WU_EXTD_TUPLE_MSB - `MGR_WU_EXTD_TUPLE_LSB +1)
`define MGR_WU_EXTD_TUPLE_RANGE             `MGR_WU_EXTD_TUPLE_MSB : `MGR_WU_EXTD_TUPLE_LSB

`define MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_MSB              `MGR_WU_EXTD_TUPLE_MSB
`define MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_LSB              `MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_MSB-(`MGR_WU_OPT_TYPE_WIDTH-1)                 
`define MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_SIZE             (`MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_MSB - `MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_LSB +1)
`define MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_RANGE             `MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_MSB : `MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_LSB

`define MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_MSB              `MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_LSB-1
`define MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_LSB              `MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_MSB-(`MGR_WU_EXTD_OPT_VALUE_WIDTH-1)
`define MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_SIZE             (`MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_MSB - `MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_LSB +1)
`define MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_RANGE             `MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_MSB : `MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_LSB


// Instruction fields
`define MGR_INST_TYPE_WIDTH               5
`define MGR_INST_TYPE_MSB                `MGR_INST_TYPE_WIDTH-1
`define MGR_INST_TYPE_LSB                 0
`define MGR_INST_TYPE_SIZE              (`MGR_INST_TYPE_MSB - `MGR_INST_TYPE_LSB +1)
`define MGR_INST_TYPE_RANGE              `MGR_INST_TYPE_MSB : `MGR_INST_TYPE_LSB

//-------------------------------------------------------------
//-------------------------------------------------------------
//-------------------------------------------------------------
// - FIXME : Must match python_typedef.vh python_desc_type
`define MGR_INST_DESC_TYPE_NOP              0
`define MGR_INST_DESC_TYPE_OP               1
`define MGR_INST_DESC_TYPE_MR               2
`define MGR_INST_DESC_TYPE_MW               3

//-------------------------------------------------------------
// - FIXME : Must match python_typedef.vh python_option_type
`define MGR_INST_OPTION_TYPE_NOP            0
`define MGR_INST_OPTION_TYPE_SRC            1
`define MGR_INST_OPTION_TYPE_TGT            2
`define MGR_INST_OPTION_TYPE_TXFER          3
`define MGR_INST_OPTION_TYPE_NUM_OF_LANES   4
`define MGR_INST_OPTION_TYPE_STOP           5
`define MGR_INST_OPTION_TYPE_SIMDOP         6
`define MGR_INST_OPTION_TYPE_MEMORY         7

//-------------------------------------------------------------
// - FIXME : Must match python_typedef.vh python_simd_type
`define MGR_INST_OPTION_SIMD_TYPE_NOP       0
`define MGR_INST_OPTION_SIMD_TYPE_RELU      1

//-------------------------------------------------------------
// - FIXME : Must match python_typedef.vh python_stOp_type
`define MGR_INST_OPTION_STOP_TYPE_NOP                                                  0
`define MGR_INST_OPTION_STOP_TYPE_STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM    1
`define MGR_INST_OPTION_STOP_TYPE_STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM      2
`define MGR_INST_OPTION_STOP_TYPE_STREAMING_OP_CNTL_OPERATION_MEM_STD_FP_MAC_TO_MEM    3

//-------------------------------------------------------------
// - FIXME : Must match python_typedef.vh python_target_type
`define MGR_INST_OPTION_TGT_TYPE_STACK_DN_ARG0   0
`define MGR_INST_OPTION_TGT_TYPE_STACK_DN_ARG1   1
`define MGR_INST_OPTION_TGT_TYPE_STACK_UP        2
`define MGR_INST_OPTION_TGT_TYPE_NOP             3


`define MGR_INST_OPTION_TGT_WIDTH        2
`define MGR_INST_OPTION_TGT_MSB          `MGR_INST_OPTION_TGT_WIDTH-1
`define MGR_INST_OPTION_TGT_LSB          0
`define MGR_INST_OPTION_TGT_SIZE         (`MGR_INST_OPTION_TGT_MSB - `MGR_INST_OPTION_TGT_LSB +1)
`define MGR_INST_OPTION_TGT_RANGE         `MGR_INST_OPTION_TGT_MSB : `MGR_INST_OPTION_TGT_LSB

//-------------------------------------------------------------
// - FIXME : Must match python_typedef.vh python_transfer_type
`define MGR_INST_OPTION_TRANSFER_TYPE_BCAST    0  
`define MGR_INST_OPTION_TRANSFER_TYPE_VECTOR   1  
`define MGR_INST_OPTION_TRANSFER_TYPE_NOP      2  

`define MGR_INST_OPTION_TRANSFER_WIDTH        2
`define MGR_INST_OPTION_TRANSFER_MSB          `MGR_INST_OPTION_TRANSFER_WIDTH-1
`define MGR_INST_OPTION_TRANSFER_LSB          0
`define MGR_INST_OPTION_TRANSFER_SIZE         (`MGR_INST_OPTION_TRANSFER_MSB - `MGR_INST_OPTION_TRANSFER_LSB +1)
`define MGR_INST_OPTION_TRANSFER_RANGE         `MGR_INST_OPTION_TRANSFER_MSB : `MGR_INST_OPTION_TRANSFER_LSB
//-------------------------------------------------------------
// - FIXME : Must match python_typedef.vh python_order_type
`define MGR_INST_OPTION_ORDER_TYPE_CWBP    0      
`define MGR_INST_OPTION_ORDER_TYPE_WCBP    1      
`define MGR_INST_OPTION_ORDER_TYPE_NOP     2      

`define MGR_INST_OPTION_ORDER_WIDTH        3
`define MGR_INST_OPTION_ORDER_MSB          `MGR_INST_OPTION_ORDER_WIDTH-1
`define MGR_INST_OPTION_ORDER_LSB          0
`define MGR_INST_OPTION_ORDER_SIZE         (`MGR_INST_OPTION_ORDER_MSB - `MGR_INST_OPTION_ORDER_LSB +1)
`define MGR_INST_OPTION_ORDER_RANGE         `MGR_INST_OPTION_ORDER_MSB : `MGR_INST_OPTION_ORDER_LSB


//---------------------------------------------------------------------------------------------------------------------
// Instruction Memory

// FIXME - need to check depth equirements (for sim, keep small)
`define MGR_INSTRUCTION_MEMORY_DEPTH   `MGR_WU_MEMORY_DEPTH 
`define MGR_INSTRUCTION_MEMORY_MSB     `MGR_INSTRUCTION_MEMORY_DEPTH-1
`define MGR_INSTRUCTION_MEMORY_LSB     0
`define MGR_INSTRUCTION_MEMORY_SIZE    (`MGR_INSTRUCTION_MEMORY_MSB - `MGR_INSTRUCTION_MEMORY_LSB +1)
`define MGR_INSTRUCTION_MEMORY_RANGE    `MGR_INSTRUCTION_MEMORY_MSB : `MGR_INSTRUCTION_MEMORY_LSB


`define MGR_INSTRUCTION_ADDRESS_WIDTH   (`CLOG2(`MGR_INSTRUCTION_MEMORY_DEPTH )) 
`define MGR_INSTRUCTION_ADDRESS_MSB     `MGR_INSTRUCTION_ADDRESS_WIDTH-1
`define MGR_INSTRUCTION_ADDRESS_LSB     0
`define MGR_INSTRUCTION_ADDRESS_SIZE    (`MGR_INSTRUCTION_ADDRESS_MSB - `MGR_INSTRUCTION_ADDRESS_LSB +1)
`define MGR_INSTRUCTION_ADDRESS_RANGE    `MGR_INSTRUCTION_ADDRESS_MSB : `MGR_INSTRUCTION_ADDRESS_LSB


`define MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_WIDTH    `COMMON_STD_INTF_CNTL_WIDTH 
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_MSB      `MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_WIDTH-1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_LSB      0
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_SIZE     (`MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_LSB +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_RANGE     `MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_LSB

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_WIDTH    `COMMON_STD_INTF_CNTL_WIDTH 
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_MSB      `MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_WIDTH-1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_LSB      `MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_MSB+1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_SIZE     (`MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_LSB +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_RANGE     `MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_LSB

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_WIDTH      `MGR_INST_TYPE_WIDTH
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_MSB      (`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_LSB+`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_WIDTH) -1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_LSB      `MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_MSB+1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_SIZE     (`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_LSB +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_RANGE     `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_LSB

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_WIDTH      `MGR_WU_OPT_TYPE_WIDTH
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_MSB      (`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_LSB+`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_WIDTH) -1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_LSB      `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_MSB+1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_SIZE     (`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_LSB +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_RANGE     `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_LSB

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_WIDTH      `MGR_WU_OPT_VALUE_WIDTH
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_MSB      (`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_LSB+`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_WIDTH) -1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_LSB      `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_MSB+1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_SIZE     (`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_LSB +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_RANGE     `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_LSB

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_WIDTH      `MGR_WU_OPT_TYPE_WIDTH
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_MSB      (`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_LSB+`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_WIDTH) -1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_LSB      `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0+1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_SIZE     (`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_LSB +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_RANGE     `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_LSB

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_WIDTH      `MGR_WU_OPT_VALUE_WIDTH
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_MSB      (`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_LSB+`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_WIDTH) -1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_LSB      `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_MSB+1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_SIZE     (`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_LSB +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_RANGE     `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_LSB

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_WIDTH      `MGR_WU_OPT_TYPE_WIDTH
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_MSB      (`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_LSB+`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_WIDTH) -1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_LSB      `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1+1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_SIZE     (`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_LSB +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_RANGE     `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_LSB

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_WIDTH      `MGR_WU_OPT_VALUE_WIDTH
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_MSB      (`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_LSB+`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_WIDTH) -1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_LSB      `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_MSB+1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_SIZE     (`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_LSB +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_RANGE     `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_LSB


`define MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_WIDTH      `MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_WIDTH     \
                                                       +`MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_WIDTH     \
                                                       +`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_WIDTH      \
                                                       +`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_WIDTH \
                                                       +`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_WIDTH  \
                                                       +`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_WIDTH \
                                                       +`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_WIDTH  \
                                                       +`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_WIDTH \
                                                       +`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_WIDTH  

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_MSB            `MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_WIDTH -1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_LSB            0
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_SIZE           (`MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_LSB +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_RANGE           `MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_LSB


//---------------------------------------------------------------------------------------------------------------------
// Storage Descriptor Memory

// FIXME - need to check depth equirements (for sim, keep small)
// This is per manager storage. The pointers will include additional bits for
// the manager ID

`define MGR_LOCAL_STORAGE_DESC_MEMORY_DEPTH   1024
`define MGR_LOCAL_STORAGE_DESC_MEMORY_MSB     `MGR_LOCAL_STORAGE_DESC_MEMORY_DEPTH-1
`define MGR_LOCAL_STORAGE_DESC_MEMORY_LSB     0
`define MGR_LOCAL_STORAGE_DESC_MEMORY_SIZE    (`MGR_LOCAL_STORAGE_DESC_MEMORY_MSB - `MGR_LOCAL_STORAGE_DESC_MEMORY_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_MEMORY_RANGE    `MGR_LOCAL_STORAGE_DESC_MEMORY_MSB : `MGR_LOCAL_STORAGE_DESC_MEMORY_LSB


`define MGR_LOCAL_STORAGE_DESC_ADDRESS_WIDTH   (`CLOG2(`MGR_LOCAL_STORAGE_DESC_MEMORY_DEPTH )) 
`define MGR_LOCAL_STORAGE_DESC_ADDRESS_MSB     `MGR_LOCAL_STORAGE_DESC_ADDRESS_WIDTH-1
`define MGR_LOCAL_STORAGE_DESC_ADDRESS_LSB     0
`define MGR_LOCAL_STORAGE_DESC_ADDRESS_SIZE    (`MGR_LOCAL_STORAGE_DESC_ADDRESS_MSB - `MGR_LOCAL_STORAGE_DESC_ADDRESS_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_ADDRESS_RANGE    `MGR_LOCAL_STORAGE_DESC_ADDRESS_MSB : `MGR_LOCAL_STORAGE_DESC_ADDRESS_LSB




// size of consequtive and jump field - FIXME : TBD
`define MGR_INST_CONS_JUMP_WIDTH        10
`define MGR_INST_CONS_JUMP_MSB          `MGR_INST_CONS_JUMP_WIDTH-1
`define MGR_INST_CONS_JUMP_LSB          0
`define MGR_INST_CONS_JUMP_SIZE         (`MGR_INST_CONS_JUMP_MSB - `MGR_INST_CONS_JUMP_LSB +1)
`define MGR_INST_CONS_JUMP_RANGE         `MGR_INST_CONS_JUMP_MSB : `MGR_INST_CONS_JUMP_LSB

// This is an array wide pointer address which has the manager id pre-pended
// Note: The pointers in the instructions are array wide pointer addresses
//
`define MGR_STORAGE_DESC_ADDRESS_WIDTH         `MGR_MGR_ID_WIDTH+`MGR_LOCAL_STORAGE_DESC_ADDRESS_WIDTH               
`define MGR_STORAGE_DESC_ADDRESS_MSB           `MGR_STORAGE_DESC_ADDRESS_WIDTH-1
`define MGR_STORAGE_DESC_ADDRESS_LSB           0
`define MGR_STORAGE_DESC_ADDRESS_SIZE          (`MGR_STORAGE_DESC_ADDRESS_MSB - `MGR_STORAGE_DESC_ADDRESS_LSB +1)
`define MGR_STORAGE_DESC_ADDRESS_RANGE          `MGR_STORAGE_DESC_ADDRESS_MSB : `MGR_STORAGE_DESC_ADDRESS_LSB

`define MGR_STORAGE_DESC_MGR_ID_FIELD_MSB      `MGR_STORAGE_DESC_ADDRESS_MSB 
`define MGR_STORAGE_DESC_MGR_ID_FIELD_LSB      `MGR_STORAGE_DESC_MGR_ID_FIELD_MSB-(`MGR_MGR_ID_WIDTH-1)
`define MGR_STORAGE_DESC_MGR_ID_FIELD_RANGE    `MGR_STORAGE_DESC_MGR_ID_FIELD_MSB : `MGR_STORAGE_DESC_MGR_ID_FIELD_LSB


// Now create aggregate memories
// FIXME: Before we can use this we need to aggregate the .dat files


`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_WIDTH    `MGR_DRAM_ADDRESS_WIDTH 
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_MSB      `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_WIDTH-1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_LSB      0
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_SIZE     (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_MSB - `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_RANGE     `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_MSB : `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_LSB

`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_WIDTH      `MGR_INST_OPTION_ORDER_WIDTH  
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_MSB      (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_LSB+`MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_WIDTH) -1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_LSB      `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_MSB+1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_SIZE     (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_MSB - `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_RANGE     `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_MSB : `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_LSB

`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_WIDTH      `MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_WIDTH 
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_MSB      (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_LSB+`MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_WIDTH) -1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_LSB      `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_MSB+1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_SIZE     (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_MSB - `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_RANGE     `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_MSB : `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_LSB


`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_WIDTH      `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_WIDTH    \
                                                       +`MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_WIDTH     \
                                                       +`MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_WIDTH    

`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_MSB            `MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_WIDTH -1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_LSB            0
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_SIZE           (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_MSB - `MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_RANGE           `MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_MSB : `MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_LSB





// Average number of consequtive/jump fields per storage descriptor
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_PER_DESC   8

`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_DEPTH   `MGR_LOCAL_STORAGE_DESC_MEMORY_DEPTH*`MGR_LOCAL_STORAGE_DESC_CONSJUMP_PER_DESC*2   // 2 ~jump,consequtive
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_MSB     `MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_DEPTH-1
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_LSB     0
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_SIZE    (`MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_MSB - `MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_RANGE    `MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_MSB : `MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_LSB


`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_WIDTH   (`CLOG2(`MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_DEPTH )) 
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_MSB     `MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_WIDTH-1
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_LSB     0
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_SIZE    (`MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_MSB - `MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_RANGE    `MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_MSB : `MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_LSB


`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_WIDTH    `MGR_INST_CONS_JUMP_WIDTH 
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_MSB      `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_WIDTH-1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_LSB      0
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_SIZE     (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_MSB - `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_RANGE     `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_MSB : `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_LSB

`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_WIDTH      `COMMON_STD_INTF_CNTL_WIDTH 
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_MSB      (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_LSB+`MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_WIDTH) -1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_LSB      `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_MSB+1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_SIZE     (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_MSB - `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_RANGE     `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_MSB : `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_LSB


`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_WIDTH       `COMMON_STD_INTF_CNTL_WIDTH   \
                                                                + `MGR_INST_CONS_JUMP_WIDTH    
                                                                

`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_MSB            `MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_WIDTH -1
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_LSB            0
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_SIZE           (`MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_MSB - `MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_RANGE           `MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_MSB : `MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_LSB















//---------------------------------------------------------------------------------------------------------------------
// DRAM Memory

`define MGR_DRAM_NUM_CHANNELS                       2
`define MGR_DRAM_NUM_BANKS                          32
`define MGR_DRAM_NUM_PAGES                          4096
`define MGR_DRAM_PAGE_SIZE                          4096
`define MGR_DRAM_NUM_WORDS_PER_PAGE                 `MGR_DRAM_PAGE_SIZE/32

// cache line size 
`define MGR_DRAM_NUM_WORDS_PER_LINE              (`MGR_DRAM_NUM_WORDS_PER_PAGE/2)
`define MGR_DRAM_NUM_LINES                       (`MGR_DRAM_NUM_WORDS_PER_PAGE/`MGR_DRAM_NUM_WORDS_PER_LINE)
//****************************************************************************************************
//****************************************************************************************************
// Note: undef MGR_DRAM_REQUEST_LT_PAGE  if an entire page is transferred during a memory access
`undef MGR_DRAM_REQUEST_LT_PAGE
`define MGR_DRAM_REQUEST_LT_PAGE
//****************************************************************************************************
//****************************************************************************************************
  

`define MGR_DRAM_NUM_CHANNELS_VECTOR_WIDTH                       `MGR_DRAM_NUM_CHANNELS
`define MGR_DRAM_NUM_CHANNELS_VECTOR_MSB                         `MGR_DRAM_NUM_CHANNELS_VECTOR_WIDTH-1
`define MGR_DRAM_NUM_CHANNELS_VECTOR_LSB                         0
`define MGR_DRAM_NUM_CHANNELS_VECTOR_SIZE                        (`MGR_DRAM_NUM_CHANNELS_VECTOR_MSB - `MGR_DRAM_NUM_CHANNELS_VECTOR_LSB +1)
`define MGR_DRAM_NUM_CHANNELS_VECTOR_RANGE                        `MGR_DRAM_NUM_CHANNELS_VECTOR_MSB : `MGR_DRAM_NUM_CHANNELS_VECTOR_LSB


//---------------------------------------------------------------------------------------------------------------------
// MMC to MRC

`define MGR_MMC_TO_MRC_INTF_WIDTH                          2048
`define MGR_MMC_TO_MRC_INTF_MSB                         `MGR_MMC_TO_MRC_INTF_WIDTH-1
`define MGR_MMC_TO_MRC_INTF_LSB                         0
`define MGR_MMC_TO_MRC_INTF_SIZE                        (`MGR_MMC_TO_MRC_INTF_MSB - `MGR_MMC_TO_MRC_INTF_LSB +1)
`define MGR_MMC_TO_MRC_INTF_RANGE                        `MGR_MMC_TO_MRC_INTF_MSB : `MGR_MMC_TO_MRC_INTF_LSB

`define MGR_MMC_TO_MRC_INTF_NUM_WORDS          `MGR_MMC_TO_MRC_INTF_WIDTH/32

`define MGR_MMC_TO_MRC_WORD_ADDRESS_WIDTH                       (`CLOG2(`MGR_MMC_TO_MRC_INTF_NUM_WORDS ))
`define MGR_MMC_TO_MRC_WORD_ADDRESS_MSB                         `MGR_MMC_TO_MRC_WORD_ADDRESS_WIDTH-1
`define MGR_MMC_TO_MRC_WORD_ADDRESS_LSB                         0
`define MGR_MMC_TO_MRC_WORD_ADDRESS_SIZE                        (`MGR_MMC_TO_MRC_WORD_ADDRESS_MSB - `MGR_MMC_TO_MRC_WORD_ADDRESS_LSB +1)
`define MGR_MMC_TO_MRC_WORD_ADDRESS_RANGE                        `MGR_MMC_TO_MRC_WORD_ADDRESS_MSB : `MGR_MMC_TO_MRC_WORD_ADDRESS_LSB

//------------------------------------------------------------------------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------------------------------------------------------------------------
// HOW MANY BITS TO ADDRESS A 64Gb MEMORY WITH 64 PORTS
//  - use byte address
//  - need to address 8GB
//  pow(2,33) = 8589934592 ~ 8G
//  we need 33 bits to address 8G e.g. 2^32 ~ 4G, + 2^31 ~ 2G + ....... + 2^0 ~ 1  ~= 8G
//  = 1

`define MGR_DRAM_CHANNEL_ADDRESS_WIDTH                       (`CLOG2(`MGR_DRAM_NUM_CHANNELS ))
`define MGR_DRAM_CHANNEL_ADDRESS_MSB                         `MGR_DRAM_CHANNEL_ADDRESS_WIDTH-1
`define MGR_DRAM_CHANNEL_ADDRESS_LSB                         0
`define MGR_DRAM_CHANNEL_ADDRESS_SIZE                        (`MGR_DRAM_CHANNEL_ADDRESS_MSB - `MGR_DRAM_CHANNEL_ADDRESS_LSB +1)
`define MGR_DRAM_CHANNEL_ADDRESS_RANGE                        `MGR_DRAM_CHANNEL_ADDRESS_MSB : `MGR_DRAM_CHANNEL_ADDRESS_LSB

`define MGR_DRAM_BANK_ADDRESS_WIDTH                       (`CLOG2(`MGR_DRAM_NUM_BANKS ))
`define MGR_DRAM_BANK_ADDRESS_MSB                         `MGR_DRAM_BANK_ADDRESS_WIDTH-1
`define MGR_DRAM_BANK_ADDRESS_LSB                         0
`define MGR_DRAM_BANK_ADDRESS_SIZE                        (`MGR_DRAM_BANK_ADDRESS_MSB - `MGR_DRAM_BANK_ADDRESS_LSB +1)
`define MGR_DRAM_BANK_ADDRESS_RANGE                        `MGR_DRAM_BANK_ADDRESS_MSB : `MGR_DRAM_BANK_ADDRESS_LSB

`define MGR_DRAM_PAGE_ADDRESS_WIDTH                      (`CLOG2(`MGR_DRAM_NUM_PAGES ))
`define MGR_DRAM_PAGE_ADDRESS_MSB                         `MGR_DRAM_PAGE_ADDRESS_WIDTH-1
`define MGR_DRAM_PAGE_ADDRESS_LSB                         0
`define MGR_DRAM_PAGE_ADDRESS_SIZE                        (`MGR_DRAM_PAGE_ADDRESS_MSB - `MGR_DRAM_PAGE_ADDRESS_LSB +1)
`define MGR_DRAM_PAGE_ADDRESS_RANGE                        `MGR_DRAM_PAGE_ADDRESS_MSB : `MGR_DRAM_PAGE_ADDRESS_LSB

`define MGR_DRAM_WORD_ADDRESS_WIDTH                       (`CLOG2(`MGR_DRAM_NUM_WORDS_PER_PAGE ))
`define MGR_DRAM_WORD_ADDRESS_MSB                         `MGR_DRAM_WORD_ADDRESS_WIDTH-1
`define MGR_DRAM_WORD_ADDRESS_LSB                         0
`define MGR_DRAM_WORD_ADDRESS_SIZE                        (`MGR_DRAM_WORD_ADDRESS_MSB - `MGR_DRAM_WORD_ADDRESS_LSB +1)
`define MGR_DRAM_WORD_ADDRESS_RANGE                        `MGR_DRAM_WORD_ADDRESS_MSB : `MGR_DRAM_WORD_ADDRESS_LSB

`ifdef  MGR_DRAM_REQUEST_LT_PAGE
  // We access a cache line for each read. We need to know which line is being accessed for the given word address in the page
  `define MGR_DRAM_LINE_ADDRESS_WIDTH                       (`CLOG2(`MGR_DRAM_NUM_LINES))
  `define MGR_DRAM_LINE_ADDRESS_MSB                         `MGR_DRAM_LINE_ADDRESS_WIDTH-1
  `define MGR_DRAM_LINE_ADDRESS_LSB                         0
  `define MGR_DRAM_LINE_ADDRESS_SIZE                        (`MGR_DRAM_LINE_ADDRESS_MSB - `MGR_DRAM_LINE_ADDRESS_LSB +1)
  `define MGR_DRAM_LINE_ADDRESS_RANGE                        `MGR_DRAM_LINE_ADDRESS_MSB : `MGR_DRAM_LINE_ADDRESS_LSB

  `define MGR_DRAM_LINE_IN_WORD_ADDRESS                    `MGR_DRAM_WORD_ADDRESS_MSB : (`MGR_DRAM_WORD_ADDRESS_MSB-(`MGR_DRAM_LINE_ADDRESS_WIDTH-1))
`endif



// DRAM has 64 interface, 2 channels,  32 banks, 4096 pages and 4096 bits per page
`define MGR_DRAM_ADDRESS_WIDTH             `MGR_MGR_ID_WIDTH+`MGR_DRAM_CHANNEL_ADDRESS_WIDTH+`MGR_DRAM_BANK_ADDRESS_WIDTH+`MGR_DRAM_PAGE_ADDRESS_WIDTH+`MGR_DRAM_WORD_ADDRESS_WIDTH+2  // byte address
`define MGR_DRAM_ADDRESS_MSB               `MGR_DRAM_ADDRESS_WIDTH-1
`define MGR_DRAM_ADDRESS_LSB               0
`define MGR_DRAM_ADDRESS_SIZE              (`MGR_DRAM_ADDRESS_MSB - `MGR_DRAM_ADDRESS_LSB +1)
`define MGR_DRAM_ADDRESS_RANGE              `MGR_DRAM_ADDRESS_MSB : `MGR_DRAM_ADDRESS_LSB

// DRAM local address width (doesnt include manager ID
`define MGR_DRAM_LOCAL_ADDRESS_WIDTH             `MGR_DRAM_CHANNEL_ADDRESS_WIDTH+`MGR_DRAM_BANK_ADDRESS_WIDTH+`MGR_DRAM_PAGE_ADDRESS_WIDTH+`MGR_DRAM_WORD_ADDRESS_WIDTH+2  // byte address
`define MGR_DRAM_LOCAL_ADDRESS_MSB               `MGR_DRAM_LOCAL_ADDRESS_WIDTH-1
`define MGR_DRAM_LOCAL_ADDRESS_LSB               0
`define MGR_DRAM_LOCAL_ADDRESS_SIZE              (`MGR_DRAM_LOCAL_ADDRESS_MSB - `MGR_DRAM_LOCAL_ADDRESS_LSB +1)
`define MGR_DRAM_LOCAL_ADDRESS_RANGE              `MGR_DRAM_LOCAL_ADDRESS_MSB : `MGR_DRAM_LOCAL_ADDRESS_LSB

// generate ranges so we can extract the fields from a given address
`define MGR_DRAM_ADDRESS_WORD_FIELD_LSB                         2  // account for byte address
`define MGR_DRAM_ADDRESS_WORD_FIELD_MSB                         `MGR_DRAM_ADDRESS_WORD_FIELD_LSB+`MGR_DRAM_WORD_ADDRESS_WIDTH-1
`define MGR_DRAM_ADDRESS_WORD_FIELD_SIZE                        (`MGR_DRAM_ADDRESS_WORD_FIELD_MSB - `MGR_DRAM_ADDRESS_WORD_FIELD_LSB +1)
`define MGR_DRAM_ADDRESS_WORD_FIELD_RANGE                        `MGR_DRAM_ADDRESS_WORD_FIELD_MSB : `MGR_DRAM_ADDRESS_WORD_FIELD_LSB

`ifdef  MGR_DRAM_REQUEST_LT_PAGE
  `define MGR_DRAM_ADDRESS_LINE_FIELD_MSB                         `MGR_DRAM_ADDRESS_WORD_FIELD_MSB
  `define MGR_DRAM_ADDRESS_LINE_FIELD_LSB                         (`MGR_DRAM_ADDRESS_LINE_FIELD_MSB-`MGR_DRAM_LINE_ADDRESS_WIDTH)+1
  `define MGR_DRAM_ADDRESS_LINE_FIELD_SIZE                        (`MGR_DRAM_ADDRESS_LINE_FIELD_MSB - `MGR_DRAM_ADDRESS_LINE_FIELD_LSB +1)
  `define MGR_DRAM_ADDRESS_LINE_FIELD_RANGE                        `MGR_DRAM_ADDRESS_LINE_FIELD_MSB : `MGR_DRAM_ADDRESS_LINE_FIELD_LSB
`endif

`define MGR_DRAM_ADDRESS_PAGE_FIELD_LSB                         `MGR_DRAM_ADDRESS_WORD_FIELD_MSB+1
`define MGR_DRAM_ADDRESS_PAGE_FIELD_MSB                         `MGR_DRAM_ADDRESS_PAGE_FIELD_LSB+`MGR_DRAM_PAGE_ADDRESS_WIDTH-1
`define MGR_DRAM_ADDRESS_PAGE_FIELD_SIZE                        (`MGR_DRAM_ADDRESS_PAGE_FIELD_MSB - `MGR_DRAM_ADDRESS_PAGE_FIELD_LSB +1)
`define MGR_DRAM_ADDRESS_PAGE_FIELD_RANGE                        `MGR_DRAM_ADDRESS_PAGE_FIELD_MSB : `MGR_DRAM_ADDRESS_PAGE_FIELD_LSB

`define MGR_DRAM_ADDRESS_BANK_FIELD_LSB                         `MGR_DRAM_ADDRESS_PAGE_FIELD_MSB+1
`define MGR_DRAM_ADDRESS_BANK_FIELD_MSB                         `MGR_DRAM_ADDRESS_BANK_FIELD_LSB+`MGR_DRAM_BANK_ADDRESS_WIDTH-1
`define MGR_DRAM_ADDRESS_BANK_FIELD_SIZE                        (`MGR_DRAM_ADDRESS_BANK_FIELD_MSB - `MGR_DRAM_ADDRESS_BANK_FIELD_LSB +1)
`define MGR_DRAM_ADDRESS_BANK_FIELD_RANGE                        `MGR_DRAM_ADDRESS_BANK_FIELD_MSB : `MGR_DRAM_ADDRESS_BANK_FIELD_LSB

`define MGR_DRAM_ADDRESS_CHAN_FIELD_LSB                         `MGR_DRAM_ADDRESS_BANK_FIELD_MSB+1
`define MGR_DRAM_ADDRESS_CHAN_FIELD_MSB                         `MGR_DRAM_ADDRESS_CHAN_FIELD_LSB+`MGR_DRAM_CHANNEL_ADDRESS_WIDTH-1
`define MGR_DRAM_ADDRESS_CHAN_FIELD_SIZE                        (`MGR_DRAM_ADDRESS_CHAN_FIELD_MSB - `MGR_DRAM_ADDRESS_CHAN_FIELD_LSB +1)
`define MGR_DRAM_ADDRESS_CHAN_FIELD_RANGE                        `MGR_DRAM_ADDRESS_CHAN_FIELD_MSB : `MGR_DRAM_ADDRESS_CHAN_FIELD_LSB

`define MGR_DRAM_ADDRESS_MGR_FIELD_LSB                         `MGR_DRAM_ADDRESS_CHAN_FIELD_MSB+1
`define MGR_DRAM_ADDRESS_MGR_FIELD_MSB                         `MGR_DRAM_ADDRESS_MGR_FIELD_LSB+`MGR_MGR_ID_WIDTH-1
`define MGR_DRAM_ADDRESS_MGR_FIELD_SIZE                        (`MGR_DRAM_ADDRESS_MGR_FIELD_MSB - `MGR_DRAM_ADDRESS_MGR_FIELD_LSB +1)
`define MGR_DRAM_ADDRESS_MGR_FIELD_RANGE                        `MGR_DRAM_ADDRESS_MGR_FIELD_MSB : `MGR_DRAM_ADDRESS_MGR_FIELD_LSB

// Field locations based on address formed from access order
// WCBP
`define MGR_DRAM_WCBP_ORDER_WORD_FIELD_LSB                         2  // account for byte address
`define MGR_DRAM_WCBP_ORDER_WORD_FIELD_MSB                         `MGR_DRAM_WCBP_ORDER_WORD_FIELD_LSB+`MGR_DRAM_WORD_ADDRESS_WIDTH-1
`define MGR_DRAM_WCBP_ORDER_WORD_FIELD_SIZE                        (`MGR_DRAM_WCBP_ORDER_WORD_FIELD_MSB - `MGR_DRAM_WCBP_ORDER_WORD_FIELD_LSB +1)
`define MGR_DRAM_WCBP_ORDER_WORD_FIELD_RANGE                        `MGR_DRAM_WCBP_ORDER_WORD_FIELD_MSB : `MGR_DRAM_WCBP_ORDER_WORD_FIELD_LSB

`define MGR_DRAM_WCBP_ORDER_CHAN_FIELD_LSB                         `MGR_DRAM_WCBP_ORDER_WORD_FIELD_MSB+1
`define MGR_DRAM_WCBP_ORDER_CHAN_FIELD_MSB                         `MGR_DRAM_WCBP_ORDER_CHAN_FIELD_LSB+`MGR_DRAM_CHANNEL_ADDRESS_WIDTH-1
`define MGR_DRAM_WCBP_ORDER_CHAN_FIELD_SIZE                        (`MGR_DRAM_WCBP_ORDER_CHAN_FIELD_MSB - `MGR_DRAM_WCBP_ORDER_CHAN_FIELD_LSB +1)
`define MGR_DRAM_WCBP_ORDER_CHAN_FIELD_RANGE                        `MGR_DRAM_WCBP_ORDER_CHAN_FIELD_MSB : `MGR_DRAM_WCBP_ORDER_CHAN_FIELD_LSB

`define MGR_DRAM_WCBP_ORDER_LINE_FIELD_LSB                         (`MGR_DRAM_WCBP_ORDER_LINE_FIELD_MSB-`MGR_DRAM_LINE_ADDRESS_WIDTH)+1
`define MGR_DRAM_WCBP_ORDER_LINE_FIELD_MSB                         `MGR_DRAM_WCBP_ORDER_WORD_FIELD_MSB
`define MGR_DRAM_WCBP_ORDER_LINE_FIELD_SIZE                        (`MGR_DRAM_WCBP_ORDER_LINE_FIELD_MSB - `MGR_DRAM_WCBP_ORDER_LINE_FIELD_LSB +1)
`define MGR_DRAM_WCBP_ORDER_LINE_FIELD_RANGE                        `MGR_DRAM_WCBP_ORDER_LINE_FIELD_MSB : `MGR_DRAM_WCBP_ORDER_LINE_FIELD_LSB

`define MGR_DRAM_WCBP_ORDER_BANK_FIELD_LSB                         `MGR_DRAM_WCBP_ORDER_CHAN_FIELD_MSB+1
`define MGR_DRAM_WCBP_ORDER_BANK_FIELD_MSB                         `MGR_DRAM_WCBP_ORDER_BANK_FIELD_LSB+`MGR_DRAM_BANK_ADDRESS_WIDTH-1
`define MGR_DRAM_WCBP_ORDER_BANK_FIELD_SIZE                        (`MGR_DRAM_WCBP_ORDER_BANK_FIELD_MSB - `MGR_DRAM_WCBP_ORDER_BANK_FIELD_LSB +1)
`define MGR_DRAM_WCBP_ORDER_BANK_FIELD_RANGE                        `MGR_DRAM_WCBP_ORDER_BANK_FIELD_MSB : `MGR_DRAM_WCBP_ORDER_BANK_FIELD_LSB

`define MGR_DRAM_WCBP_ORDER_PAGE_FIELD_LSB                         `MGR_DRAM_WCBP_ORDER_BANK_FIELD_MSB+1
`define MGR_DRAM_WCBP_ORDER_PAGE_FIELD_MSB                         `MGR_DRAM_WCBP_ORDER_PAGE_FIELD_LSB+`MGR_DRAM_PAGE_ADDRESS_WIDTH-1
`define MGR_DRAM_WCBP_ORDER_PAGE_FIELD_SIZE                        (`MGR_DRAM_WCBP_ORDER_PAGE_FIELD_MSB - `MGR_DRAM_WCBP_ORDER_PAGE_FIELD_LSB +1)
`define MGR_DRAM_WCBP_ORDER_PAGE_FIELD_RANGE                        `MGR_DRAM_WCBP_ORDER_PAGE_FIELD_MSB : `MGR_DRAM_WCBP_ORDER_PAGE_FIELD_LSB


// CWBP
`define MGR_DRAM_CWBP_ORDER_CHAN_FIELD_LSB                         2  // account for byte address
`define MGR_DRAM_CWBP_ORDER_CHAN_FIELD_MSB                         `MGR_DRAM_CWBP_ORDER_CHAN_FIELD_LSB+`MGR_DRAM_CHANNEL_ADDRESS_WIDTH-1
`define MGR_DRAM_CWBP_ORDER_CHAN_FIELD_SIZE                        (`MGR_DRAM_CWBP_ORDER_CHAN_FIELD_MSB - `MGR_DRAM_CWBP_ORDER_CHAN_FIELD_LSB +1)
`define MGR_DRAM_CWBP_ORDER_CHAN_FIELD_RANGE                        `MGR_DRAM_CWBP_ORDER_CHAN_FIELD_MSB : `MGR_DRAM_CWBP_ORDER_CHAN_FIELD_LSB

`define MGR_DRAM_CWBP_ORDER_WORD_FIELD_LSB                         `MGR_DRAM_CWBP_ORDER_CHAN_FIELD_MSB+1
`define MGR_DRAM_CWBP_ORDER_WORD_FIELD_MSB                         `MGR_DRAM_CWBP_ORDER_WORD_FIELD_LSB+`MGR_DRAM_WORD_ADDRESS_WIDTH-1
`define MGR_DRAM_CWBP_ORDER_WORD_FIELD_SIZE                        (`MGR_DRAM_CWBP_ORDER_WORD_FIELD_MSB - `MGR_DRAM_CWBP_ORDER_WORD_FIELD_LSB +1)
`define MGR_DRAM_CWBP_ORDER_WORD_FIELD_RANGE                        `MGR_DRAM_CWBP_ORDER_WORD_FIELD_MSB : `MGR_DRAM_CWBP_ORDER_WORD_FIELD_LSB

`define MGR_DRAM_CWBP_ORDER_LINE_FIELD_LSB                         (`MGR_DRAM_CWBP_ORDER_LINE_FIELD_MSB-`MGR_DRAM_LINE_ADDRESS_WIDTH)+1
`define MGR_DRAM_CWBP_ORDER_LINE_FIELD_MSB                         `MGR_DRAM_CWBP_ORDER_WORD_FIELD_MSB
`define MGR_DRAM_CWBP_ORDER_LINE_FIELD_SIZE                        (`MGR_DRAM_CWBP_ORDER_LINE_FIELD_MSB - `MGR_DRAM_CWBP_ORDER_LINE_FIELD_LSB +1)
`define MGR_DRAM_CWBP_ORDER_LINE_FIELD_RANGE                        `MGR_DRAM_CWBP_ORDER_LINE_FIELD_MSB : `MGR_DRAM_CWBP_ORDER_LINE_FIELD_LSB

`define MGR_DRAM_CWBP_ORDER_BANK_FIELD_LSB                         `MGR_DRAM_CWBP_ORDER_WORD_FIELD_MSB+1
`define MGR_DRAM_CWBP_ORDER_BANK_FIELD_MSB                         `MGR_DRAM_CWBP_ORDER_BANK_FIELD_LSB+`MGR_DRAM_BANK_ADDRESS_WIDTH-1
`define MGR_DRAM_CWBP_ORDER_BANK_FIELD_SIZE                        (`MGR_DRAM_CWBP_ORDER_BANK_FIELD_MSB - `MGR_DRAM_CWBP_ORDER_BANK_FIELD_LSB +1)
`define MGR_DRAM_CWBP_ORDER_BANK_FIELD_RANGE                        `MGR_DRAM_CWBP_ORDER_BANK_FIELD_MSB : `MGR_DRAM_CWBP_ORDER_BANK_FIELD_LSB

`define MGR_DRAM_CWBP_ORDER_PAGE_FIELD_LSB                         `MGR_DRAM_CWBP_ORDER_BANK_FIELD_MSB+1
`define MGR_DRAM_CWBP_ORDER_PAGE_FIELD_MSB                         `MGR_DRAM_CWBP_ORDER_PAGE_FIELD_LSB+`MGR_DRAM_PAGE_ADDRESS_WIDTH-1
`define MGR_DRAM_CWBP_ORDER_PAGE_FIELD_SIZE                        (`MGR_DRAM_CWBP_ORDER_PAGE_FIELD_MSB - `MGR_DRAM_CWBP_ORDER_PAGE_FIELD_LSB +1)
`define MGR_DRAM_CWBP_ORDER_PAGE_FIELD_RANGE                        `MGR_DRAM_CWBP_ORDER_PAGE_FIELD_MSB : `MGR_DRAM_CWBP_ORDER_PAGE_FIELD_LSB

//------------------------------------------------------------------------------------------------------------------------
// The memory requestor will always open the next channel/bank/page based on the current address
// If a memory request provides an entire page, then to determine whether we
// need a request, just form an adrress based on page/bank/channel and increment 
// If a memry request is a partial page (line), then form an address based on PBLC or PBCL
//
// 1) Line same size as page, so only increment page/bank/channel
// PBC
`define MGR_DRAM_PBC_CHAN_FIELD_WIDTH       `MGR_DRAM_CHANNEL_ADDRESS_WIDTH
`define MGR_DRAM_PBC_CHAN_FIELD_LSB         0
`define MGR_DRAM_PBC_CHAN_FIELD_MSB         `MGR_DRAM_PBC_CHAN_FIELD_LSB+`MGR_DRAM_PBC_CHAN_FIELD_WIDTH -1
`define MGR_DRAM_PBC_CHAN_FIELD_SIZE        (`MGR_DRAM_PBC_CHAN_FIELD_MSB - `MGR_DRAM_PBC_CHAN_FIELD_LSB +1)
`define MGR_DRAM_PBC_CHAN_FIELD_RANGE        `MGR_DRAM_PBC_CHAN_FIELD_MSB : `MGR_DRAM_PBC_CHAN_FIELD_LSB

`define MGR_DRAM_PBC_BANK_FIELD_WIDTH       `MGR_DRAM_BANK_ADDRESS_WIDTH
`define MGR_DRAM_PBC_BANK_FIELD_LSB         `MGR_DRAM_PBC_CHAN_FIELD_MSB+1
`define MGR_DRAM_PBC_BANK_FIELD_MSB         `MGR_DRAM_PBC_BANK_FIELD_LSB+`MGR_DRAM_PBC_BANK_FIELD_WIDTH -1
`define MGR_DRAM_PBC_BANK_FIELD_SIZE        (`MGR_DRAM_PBC_BANK_FIELD_MSB - `MGR_DRAM_PBC_BANK_FIELD_LSB +1)
`define MGR_DRAM_PBC_BANK_FIELD_RANGE        `MGR_DRAM_PBC_BANK_FIELD_MSB : `MGR_DRAM_PBC_BANK_FIELD_LSB

`define MGR_DRAM_PBC_PAGE_FIELD_WIDTH       `MGR_DRAM_PAGE_ADDRESS_WIDTH
`define MGR_DRAM_PBC_PAGE_FIELD_LSB         `MGR_DRAM_PBC_BANK_FIELD_MSB+1
`define MGR_DRAM_PBC_PAGE_FIELD_MSB         `MGR_DRAM_PBC_PAGE_FIELD_LSB+`MGR_DRAM_PBC_PAGE_FIELD_WIDTH -1
`define MGR_DRAM_PBC_PAGE_FIELD_SIZE        (`MGR_DRAM_PBC_PAGE_FIELD_MSB - `MGR_DRAM_PBC_PAGE_FIELD_LSB +1)
`define MGR_DRAM_PBC_PAGE_FIELD_RANGE        `MGR_DRAM_PBC_PAGE_FIELD_MSB : `MGR_DRAM_PBC_PAGE_FIELD_LSB

`define MGR_DRAM_PBC_WIDTH                   `MGR_DRAM_PBC_PAGE_FIELD_WIDTH      \
                                            +`MGR_DRAM_PBC_BANK_FIELD_WIDTH      \
                                            +`MGR_DRAM_PBC_CHAN_FIELD_WIDTH 
                                            
`define MGR_DRAM_PBC_MSB            `MGR_DRAM_PBC_WIDTH -1
`define MGR_DRAM_PBC_LSB            0
`define MGR_DRAM_PBC_SIZE           (`MGR_DRAM_PBC_MSB - `MGR_DRAM_PBC_LSB +1)
`define MGR_DRAM_PBC_RANGE           `MGR_DRAM_PBC_MSB : `MGR_DRAM_PBC_LSB



// 2) Line smaller than page, so increment either page/bank/channel/line or page/bank/line/channel
`ifdef  MGR_DRAM_REQUEST_LT_PAGE

  //----------------------------------------------------------------------------------------------------
  // PBCL
  `define MGR_DRAM_PBCL_LINE_FIELD_WIDTH       `MGR_DRAM_LINE_ADDRESS_WIDTH 
  `define MGR_DRAM_PBCL_LINE_FIELD_LSB         0
  `define MGR_DRAM_PBCL_LINE_FIELD_MSB         `MGR_DRAM_PBCL_LINE_FIELD_LSB+`MGR_DRAM_PBCL_LINE_FIELD_WIDTH -1
  `define MGR_DRAM_PBCL_LINE_FIELD_SIZE        (`MGR_DRAM_PBCL_LINE_FIELD_MSB - `MGR_DRAM_PBCL_LINE_FIELD_LSB +1)
  `define MGR_DRAM_PBCL_LINE_FIELD_RANGE        `MGR_DRAM_PBCL_LINE_FIELD_MSB : `MGR_DRAM_PBCL_LINE_FIELD_LSB

  `define MGR_DRAM_PBCL_CHAN_FIELD_WIDTH       `MGR_DRAM_CHANNEL_ADDRESS_WIDTH
  `define MGR_DRAM_PBCL_CHAN_FIELD_LSB         `MGR_DRAM_PBCL_LINE_FIELD_MSB+1
  `define MGR_DRAM_PBCL_CHAN_FIELD_MSB         `MGR_DRAM_PBCL_CHAN_FIELD_LSB+`MGR_DRAM_PBCL_CHAN_FIELD_WIDTH -1
  `define MGR_DRAM_PBCL_CHAN_FIELD_SIZE        (`MGR_DRAM_PBCL_CHAN_FIELD_MSB - `MGR_DRAM_PBCL_CHAN_FIELD_LSB +1)
  `define MGR_DRAM_PBCL_CHAN_FIELD_RANGE        `MGR_DRAM_PBCL_CHAN_FIELD_MSB : `MGR_DRAM_PBCL_CHAN_FIELD_LSB
  
  `define MGR_DRAM_PBCL_BANK_FIELD_WIDTH       `MGR_DRAM_BANK_ADDRESS_WIDTH
  `define MGR_DRAM_PBCL_BANK_FIELD_LSB         `MGR_DRAM_PBCL_CHAN_FIELD_MSB+1
  `define MGR_DRAM_PBCL_BANK_FIELD_MSB         `MGR_DRAM_PBCL_BANK_FIELD_LSB+`MGR_DRAM_PBCL_BANK_FIELD_WIDTH -1
  `define MGR_DRAM_PBCL_BANK_FIELD_SIZE        (`MGR_DRAM_PBCL_BANK_FIELD_MSB - `MGR_DRAM_PBCL_BANK_FIELD_LSB +1)
  `define MGR_DRAM_PBCL_BANK_FIELD_RANGE        `MGR_DRAM_PBCL_BANK_FIELD_MSB : `MGR_DRAM_PBCL_BANK_FIELD_LSB
  
  `define MGR_DRAM_PBCL_PAGE_FIELD_WIDTH       `MGR_DRAM_PAGE_ADDRESS_WIDTH
  `define MGR_DRAM_PBCL_PAGE_FIELD_LSB         `MGR_DRAM_PBCL_BANK_FIELD_MSB+1
  `define MGR_DRAM_PBCL_PAGE_FIELD_MSB         `MGR_DRAM_PBCL_PAGE_FIELD_LSB+`MGR_DRAM_PBCL_PAGE_FIELD_WIDTH -1
  `define MGR_DRAM_PBCL_PAGE_FIELD_SIZE        (`MGR_DRAM_PBCL_PAGE_FIELD_MSB - `MGR_DRAM_PBCL_PAGE_FIELD_LSB +1)
  `define MGR_DRAM_PBCL_PAGE_FIELD_RANGE        `MGR_DRAM_PBCL_PAGE_FIELD_MSB : `MGR_DRAM_PBCL_PAGE_FIELD_LSB
  
  `define MGR_DRAM_PBCL_WIDTH                   `MGR_DRAM_PBCL_PAGE_FIELD_WIDTH      \
                                               +`MGR_DRAM_PBCL_BANK_FIELD_WIDTH      \
                                               +`MGR_DRAM_PBCL_CHAN_FIELD_WIDTH      \
                                               +`MGR_DRAM_PBCL_LINE_FIELD_WIDTH       
  
  
  `define MGR_DRAM_PBCL_MSB            `MGR_DRAM_PBCL_WIDTH -1
  `define MGR_DRAM_PBCL_LSB            0
  `define MGR_DRAM_PBCL_SIZE           (`MGR_DRAM_PBCL_MSB - `MGR_DRAM_PBCL_LSB +1)
  `define MGR_DRAM_PBCL_RANGE           `MGR_DRAM_PBCL_MSB : `MGR_DRAM_PBCL_LSB

  //----------------------------------------------------------------------------------------------------
  // PBLC
  `define MGR_DRAM_PBLC_CHAN_FIELD_WIDTH       `MGR_DRAM_CHANNEL_ADDRESS_WIDTH
  `define MGR_DRAM_PBLC_CHAN_FIELD_LSB         0
  `define MGR_DRAM_PBLC_CHAN_FIELD_MSB         `MGR_DRAM_PBLC_CHAN_FIELD_LSB+`MGR_DRAM_PBLC_CHAN_FIELD_WIDTH -1
  `define MGR_DRAM_PBLC_CHAN_FIELD_SIZE        (`MGR_DRAM_PBLC_CHAN_FIELD_MSB - `MGR_DRAM_PBLC_CHAN_FIELD_LSB +1)
  `define MGR_DRAM_PBLC_CHAN_FIELD_RANGE        `MGR_DRAM_PBLC_CHAN_FIELD_MSB : `MGR_DRAM_PBLC_CHAN_FIELD_LSB
  
  `define MGR_DRAM_PBLC_LINE_FIELD_WIDTH       `MGR_DRAM_LINE_ADDRESS_WIDTH 
  `define MGR_DRAM_PBLC_LINE_FIELD_LSB         `MGR_DRAM_PBLC_CHAN_FIELD_MSB+1
  `define MGR_DRAM_PBLC_LINE_FIELD_MSB         `MGR_DRAM_PBLC_LINE_FIELD_LSB+`MGR_DRAM_PBLC_LINE_FIELD_WIDTH -1
  `define MGR_DRAM_PBLC_LINE_FIELD_SIZE        (`MGR_DRAM_PBLC_LINE_FIELD_MSB - `MGR_DRAM_PBLC_LINE_FIELD_LSB +1)
  `define MGR_DRAM_PBLC_LINE_FIELD_RANGE        `MGR_DRAM_PBLC_LINE_FIELD_MSB : `MGR_DRAM_PBLC_LINE_FIELD_LSB

  `define MGR_DRAM_PBLC_BANK_FIELD_WIDTH       `MGR_DRAM_BANK_ADDRESS_WIDTH
  `define MGR_DRAM_PBLC_BANK_FIELD_LSB         `MGR_DRAM_PBLC_LINE_FIELD_MSB+1
  `define MGR_DRAM_PBLC_BANK_FIELD_MSB         `MGR_DRAM_PBLC_BANK_FIELD_LSB+`MGR_DRAM_PBLC_BANK_FIELD_WIDTH -1
  `define MGR_DRAM_PBLC_BANK_FIELD_SIZE        (`MGR_DRAM_PBLC_BANK_FIELD_MSB - `MGR_DRAM_PBLC_BANK_FIELD_LSB +1)
  `define MGR_DRAM_PBLC_BANK_FIELD_RANGE        `MGR_DRAM_PBLC_BANK_FIELD_MSB : `MGR_DRAM_PBLC_BANK_FIELD_LSB
  
  `define MGR_DRAM_PBLC_PAGE_FIELD_WIDTH       `MGR_DRAM_PAGE_ADDRESS_WIDTH
  `define MGR_DRAM_PBLC_PAGE_FIELD_LSB         `MGR_DRAM_PBLC_BANK_FIELD_MSB+1
  `define MGR_DRAM_PBLC_PAGE_FIELD_MSB         `MGR_DRAM_PBLC_PAGE_FIELD_LSB+`MGR_DRAM_PBLC_PAGE_FIELD_WIDTH -1
  `define MGR_DRAM_PBLC_PAGE_FIELD_SIZE        (`MGR_DRAM_PBLC_PAGE_FIELD_MSB - `MGR_DRAM_PBLC_PAGE_FIELD_LSB +1)
  `define MGR_DRAM_PBLC_PAGE_FIELD_RANGE        `MGR_DRAM_PBLC_PAGE_FIELD_MSB : `MGR_DRAM_PBLC_PAGE_FIELD_LSB
  
  `define MGR_DRAM_PBLC_WIDTH                   `MGR_DRAM_PBLC_PAGE_FIELD_WIDTH      \
                                               +`MGR_DRAM_PBLC_BANK_FIELD_WIDTH      \
                                               +`MGR_DRAM_PBLC_CHAN_FIELD_WIDTH      \
                                               +`MGR_DRAM_PBLC_LINE_FIELD_WIDTH       
  
  
  `define MGR_DRAM_PBLC_MSB            `MGR_DRAM_PBLC_WIDTH -1
  `define MGR_DRAM_PBLC_LSB            0
  `define MGR_DRAM_PBLC_SIZE           (`MGR_DRAM_PBLC_MSB - `MGR_DRAM_PBLC_LSB +1)
  `define MGR_DRAM_PBLC_RANGE           `MGR_DRAM_PBLC_MSB : `MGR_DRAM_PBLC_LSB


`endif


//---------------------------------------------------------------------------------------------------------------------
// NoC

`define MGR_NOC_INTERNAL_DATA_WIDTH        `MGR_ARRAY_NOC_INTERNAL_DATA_WIDTH
`define MGR_NOC_INTERNAL_DATA_MSB          `MGR_NOC_INTERNAL_DATA_WIDTH-1
`define MGR_NOC_INTERNAL_DATA_LSB          0
`define MGR_NOC_INTERNAL_DATA_RANGE        `MGR_NOC_INTERNAL_DATA_MSB : `MGR_NOC_INTERNAL_DATA_LSB

`define MGR_NOC_EXTERNAL_DATA_WIDTH        `MGR_ARRAY_NOC_EXTERNAL_DATA_WIDTH 
`define MGR_NOC_EXTERNAL_DATA_MSB          `MGR_NOC_EXTERNAL_DATA_WIDTH-1
`define MGR_NOC_EXTERNAL_DATA_LSB          0
`define MGR_NOC_EXTERNAL_DATA_RANGE        `MGR_NOC_EXTERNAL_DATA_MSB : `MGR_NOC_EXTERNAL_DATA_LSB


//---------------------------------------------------------------------------------------------------------------------



`endif
