
  // General control and status                                                  
  input                                         sys__pe0__allSynchronized     ;
  output                                        pe0__sys__thisSynchronized    ;
  output                                        pe0__sys__ready               ;
  output                                        pe0__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe1__allSynchronized     ;
  output                                        pe1__sys__thisSynchronized    ;
  output                                        pe1__sys__ready               ;
  output                                        pe1__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe2__allSynchronized     ;
  output                                        pe2__sys__thisSynchronized    ;
  output                                        pe2__sys__ready               ;
  output                                        pe2__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe3__allSynchronized     ;
  output                                        pe3__sys__thisSynchronized    ;
  output                                        pe3__sys__ready               ;
  output                                        pe3__sys__complete            ;