
  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe0__allSynchronized    ( DownstreamStackBusOOB[0].cb_test.sys__pe__allSynchronized   ), 
        .pe0__sys__thisSynchronized   ( DownstreamStackBusOOB[0].pe__sys__thisSynchronized          ), 
        .pe0__sys__ready              ( DownstreamStackBusOOB[0].pe__sys__ready                     ), 
        .pe0__sys__complete           ( DownstreamStackBusOOB[0].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe1__allSynchronized    ( DownstreamStackBusOOB[1].cb_test.sys__pe__allSynchronized   ), 
        .pe1__sys__thisSynchronized   ( DownstreamStackBusOOB[1].pe__sys__thisSynchronized          ), 
        .pe1__sys__ready              ( DownstreamStackBusOOB[1].pe__sys__ready                     ), 
        .pe1__sys__complete           ( DownstreamStackBusOOB[1].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe2__allSynchronized    ( DownstreamStackBusOOB[2].cb_test.sys__pe__allSynchronized   ), 
        .pe2__sys__thisSynchronized   ( DownstreamStackBusOOB[2].pe__sys__thisSynchronized          ), 
        .pe2__sys__ready              ( DownstreamStackBusOOB[2].pe__sys__ready                     ), 
        .pe2__sys__complete           ( DownstreamStackBusOOB[2].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe3__allSynchronized    ( DownstreamStackBusOOB[3].cb_test.sys__pe__allSynchronized   ), 
        .pe3__sys__thisSynchronized   ( DownstreamStackBusOOB[3].pe__sys__thisSynchronized          ), 
        .pe3__sys__ready              ( DownstreamStackBusOOB[3].pe__sys__ready                     ), 
        .pe3__sys__complete           ( DownstreamStackBusOOB[3].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe4__allSynchronized    ( DownstreamStackBusOOB[4].cb_test.sys__pe__allSynchronized   ), 
        .pe4__sys__thisSynchronized   ( DownstreamStackBusOOB[4].pe__sys__thisSynchronized          ), 
        .pe4__sys__ready              ( DownstreamStackBusOOB[4].pe__sys__ready                     ), 
        .pe4__sys__complete           ( DownstreamStackBusOOB[4].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe5__allSynchronized    ( DownstreamStackBusOOB[5].cb_test.sys__pe__allSynchronized   ), 
        .pe5__sys__thisSynchronized   ( DownstreamStackBusOOB[5].pe__sys__thisSynchronized          ), 
        .pe5__sys__ready              ( DownstreamStackBusOOB[5].pe__sys__ready                     ), 
        .pe5__sys__complete           ( DownstreamStackBusOOB[5].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe6__allSynchronized    ( DownstreamStackBusOOB[6].cb_test.sys__pe__allSynchronized   ), 
        .pe6__sys__thisSynchronized   ( DownstreamStackBusOOB[6].pe__sys__thisSynchronized          ), 
        .pe6__sys__ready              ( DownstreamStackBusOOB[6].pe__sys__ready                     ), 
        .pe6__sys__complete           ( DownstreamStackBusOOB[6].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe7__allSynchronized    ( DownstreamStackBusOOB[7].cb_test.sys__pe__allSynchronized   ), 
        .pe7__sys__thisSynchronized   ( DownstreamStackBusOOB[7].pe__sys__thisSynchronized          ), 
        .pe7__sys__ready              ( DownstreamStackBusOOB[7].pe__sys__ready                     ), 
        .pe7__sys__complete           ( DownstreamStackBusOOB[7].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe8__allSynchronized    ( DownstreamStackBusOOB[8].cb_test.sys__pe__allSynchronized   ), 
        .pe8__sys__thisSynchronized   ( DownstreamStackBusOOB[8].pe__sys__thisSynchronized          ), 
        .pe8__sys__ready              ( DownstreamStackBusOOB[8].pe__sys__ready                     ), 
        .pe8__sys__complete           ( DownstreamStackBusOOB[8].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe9__allSynchronized    ( DownstreamStackBusOOB[9].cb_test.sys__pe__allSynchronized   ), 
        .pe9__sys__thisSynchronized   ( DownstreamStackBusOOB[9].pe__sys__thisSynchronized          ), 
        .pe9__sys__ready              ( DownstreamStackBusOOB[9].pe__sys__ready                     ), 
        .pe9__sys__complete           ( DownstreamStackBusOOB[9].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe10__allSynchronized    ( DownstreamStackBusOOB[10].cb_test.sys__pe__allSynchronized   ), 
        .pe10__sys__thisSynchronized   ( DownstreamStackBusOOB[10].pe__sys__thisSynchronized          ), 
        .pe10__sys__ready              ( DownstreamStackBusOOB[10].pe__sys__ready                     ), 
        .pe10__sys__complete           ( DownstreamStackBusOOB[10].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe11__allSynchronized    ( DownstreamStackBusOOB[11].cb_test.sys__pe__allSynchronized   ), 
        .pe11__sys__thisSynchronized   ( DownstreamStackBusOOB[11].pe__sys__thisSynchronized          ), 
        .pe11__sys__ready              ( DownstreamStackBusOOB[11].pe__sys__ready                     ), 
        .pe11__sys__complete           ( DownstreamStackBusOOB[11].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe12__allSynchronized    ( DownstreamStackBusOOB[12].cb_test.sys__pe__allSynchronized   ), 
        .pe12__sys__thisSynchronized   ( DownstreamStackBusOOB[12].pe__sys__thisSynchronized          ), 
        .pe12__sys__ready              ( DownstreamStackBusOOB[12].pe__sys__ready                     ), 
        .pe12__sys__complete           ( DownstreamStackBusOOB[12].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe13__allSynchronized    ( DownstreamStackBusOOB[13].cb_test.sys__pe__allSynchronized   ), 
        .pe13__sys__thisSynchronized   ( DownstreamStackBusOOB[13].pe__sys__thisSynchronized          ), 
        .pe13__sys__ready              ( DownstreamStackBusOOB[13].pe__sys__ready                     ), 
        .pe13__sys__complete           ( DownstreamStackBusOOB[13].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe14__allSynchronized    ( DownstreamStackBusOOB[14].cb_test.sys__pe__allSynchronized   ), 
        .pe14__sys__thisSynchronized   ( DownstreamStackBusOOB[14].pe__sys__thisSynchronized          ), 
        .pe14__sys__ready              ( DownstreamStackBusOOB[14].pe__sys__ready                     ), 
        .pe14__sys__complete           ( DownstreamStackBusOOB[14].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe15__allSynchronized    ( DownstreamStackBusOOB[15].cb_test.sys__pe__allSynchronized   ), 
        .pe15__sys__thisSynchronized   ( DownstreamStackBusOOB[15].pe__sys__thisSynchronized          ), 
        .pe15__sys__ready              ( DownstreamStackBusOOB[15].pe__sys__ready                     ), 
        .pe15__sys__complete           ( DownstreamStackBusOOB[15].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe16__allSynchronized    ( DownstreamStackBusOOB[16].cb_test.sys__pe__allSynchronized   ), 
        .pe16__sys__thisSynchronized   ( DownstreamStackBusOOB[16].pe__sys__thisSynchronized          ), 
        .pe16__sys__ready              ( DownstreamStackBusOOB[16].pe__sys__ready                     ), 
        .pe16__sys__complete           ( DownstreamStackBusOOB[16].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe17__allSynchronized    ( DownstreamStackBusOOB[17].cb_test.sys__pe__allSynchronized   ), 
        .pe17__sys__thisSynchronized   ( DownstreamStackBusOOB[17].pe__sys__thisSynchronized          ), 
        .pe17__sys__ready              ( DownstreamStackBusOOB[17].pe__sys__ready                     ), 
        .pe17__sys__complete           ( DownstreamStackBusOOB[17].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe18__allSynchronized    ( DownstreamStackBusOOB[18].cb_test.sys__pe__allSynchronized   ), 
        .pe18__sys__thisSynchronized   ( DownstreamStackBusOOB[18].pe__sys__thisSynchronized          ), 
        .pe18__sys__ready              ( DownstreamStackBusOOB[18].pe__sys__ready                     ), 
        .pe18__sys__complete           ( DownstreamStackBusOOB[18].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe19__allSynchronized    ( DownstreamStackBusOOB[19].cb_test.sys__pe__allSynchronized   ), 
        .pe19__sys__thisSynchronized   ( DownstreamStackBusOOB[19].pe__sys__thisSynchronized          ), 
        .pe19__sys__ready              ( DownstreamStackBusOOB[19].pe__sys__ready                     ), 
        .pe19__sys__complete           ( DownstreamStackBusOOB[19].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe20__allSynchronized    ( DownstreamStackBusOOB[20].cb_test.sys__pe__allSynchronized   ), 
        .pe20__sys__thisSynchronized   ( DownstreamStackBusOOB[20].pe__sys__thisSynchronized          ), 
        .pe20__sys__ready              ( DownstreamStackBusOOB[20].pe__sys__ready                     ), 
        .pe20__sys__complete           ( DownstreamStackBusOOB[20].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe21__allSynchronized    ( DownstreamStackBusOOB[21].cb_test.sys__pe__allSynchronized   ), 
        .pe21__sys__thisSynchronized   ( DownstreamStackBusOOB[21].pe__sys__thisSynchronized          ), 
        .pe21__sys__ready              ( DownstreamStackBusOOB[21].pe__sys__ready                     ), 
        .pe21__sys__complete           ( DownstreamStackBusOOB[21].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe22__allSynchronized    ( DownstreamStackBusOOB[22].cb_test.sys__pe__allSynchronized   ), 
        .pe22__sys__thisSynchronized   ( DownstreamStackBusOOB[22].pe__sys__thisSynchronized          ), 
        .pe22__sys__ready              ( DownstreamStackBusOOB[22].pe__sys__ready                     ), 
        .pe22__sys__complete           ( DownstreamStackBusOOB[22].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe23__allSynchronized    ( DownstreamStackBusOOB[23].cb_test.sys__pe__allSynchronized   ), 
        .pe23__sys__thisSynchronized   ( DownstreamStackBusOOB[23].pe__sys__thisSynchronized          ), 
        .pe23__sys__ready              ( DownstreamStackBusOOB[23].pe__sys__ready                     ), 
        .pe23__sys__complete           ( DownstreamStackBusOOB[23].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe24__allSynchronized    ( DownstreamStackBusOOB[24].cb_test.sys__pe__allSynchronized   ), 
        .pe24__sys__thisSynchronized   ( DownstreamStackBusOOB[24].pe__sys__thisSynchronized          ), 
        .pe24__sys__ready              ( DownstreamStackBusOOB[24].pe__sys__ready                     ), 
        .pe24__sys__complete           ( DownstreamStackBusOOB[24].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe25__allSynchronized    ( DownstreamStackBusOOB[25].cb_test.sys__pe__allSynchronized   ), 
        .pe25__sys__thisSynchronized   ( DownstreamStackBusOOB[25].pe__sys__thisSynchronized          ), 
        .pe25__sys__ready              ( DownstreamStackBusOOB[25].pe__sys__ready                     ), 
        .pe25__sys__complete           ( DownstreamStackBusOOB[25].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe26__allSynchronized    ( DownstreamStackBusOOB[26].cb_test.sys__pe__allSynchronized   ), 
        .pe26__sys__thisSynchronized   ( DownstreamStackBusOOB[26].pe__sys__thisSynchronized          ), 
        .pe26__sys__ready              ( DownstreamStackBusOOB[26].pe__sys__ready                     ), 
        .pe26__sys__complete           ( DownstreamStackBusOOB[26].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe27__allSynchronized    ( DownstreamStackBusOOB[27].cb_test.sys__pe__allSynchronized   ), 
        .pe27__sys__thisSynchronized   ( DownstreamStackBusOOB[27].pe__sys__thisSynchronized          ), 
        .pe27__sys__ready              ( DownstreamStackBusOOB[27].pe__sys__ready                     ), 
        .pe27__sys__complete           ( DownstreamStackBusOOB[27].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe28__allSynchronized    ( DownstreamStackBusOOB[28].cb_test.sys__pe__allSynchronized   ), 
        .pe28__sys__thisSynchronized   ( DownstreamStackBusOOB[28].pe__sys__thisSynchronized          ), 
        .pe28__sys__ready              ( DownstreamStackBusOOB[28].pe__sys__ready                     ), 
        .pe28__sys__complete           ( DownstreamStackBusOOB[28].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe29__allSynchronized    ( DownstreamStackBusOOB[29].cb_test.sys__pe__allSynchronized   ), 
        .pe29__sys__thisSynchronized   ( DownstreamStackBusOOB[29].pe__sys__thisSynchronized          ), 
        .pe29__sys__ready              ( DownstreamStackBusOOB[29].pe__sys__ready                     ), 
        .pe29__sys__complete           ( DownstreamStackBusOOB[29].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe30__allSynchronized    ( DownstreamStackBusOOB[30].cb_test.sys__pe__allSynchronized   ), 
        .pe30__sys__thisSynchronized   ( DownstreamStackBusOOB[30].pe__sys__thisSynchronized          ), 
        .pe30__sys__ready              ( DownstreamStackBusOOB[30].pe__sys__ready                     ), 
        .pe30__sys__complete           ( DownstreamStackBusOOB[30].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe31__allSynchronized    ( DownstreamStackBusOOB[31].cb_test.sys__pe__allSynchronized   ), 
        .pe31__sys__thisSynchronized   ( DownstreamStackBusOOB[31].pe__sys__thisSynchronized          ), 
        .pe31__sys__ready              ( DownstreamStackBusOOB[31].pe__sys__ready                     ), 
        .pe31__sys__complete           ( DownstreamStackBusOOB[31].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe32__allSynchronized    ( DownstreamStackBusOOB[32].cb_test.sys__pe__allSynchronized   ), 
        .pe32__sys__thisSynchronized   ( DownstreamStackBusOOB[32].pe__sys__thisSynchronized          ), 
        .pe32__sys__ready              ( DownstreamStackBusOOB[32].pe__sys__ready                     ), 
        .pe32__sys__complete           ( DownstreamStackBusOOB[32].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe33__allSynchronized    ( DownstreamStackBusOOB[33].cb_test.sys__pe__allSynchronized   ), 
        .pe33__sys__thisSynchronized   ( DownstreamStackBusOOB[33].pe__sys__thisSynchronized          ), 
        .pe33__sys__ready              ( DownstreamStackBusOOB[33].pe__sys__ready                     ), 
        .pe33__sys__complete           ( DownstreamStackBusOOB[33].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe34__allSynchronized    ( DownstreamStackBusOOB[34].cb_test.sys__pe__allSynchronized   ), 
        .pe34__sys__thisSynchronized   ( DownstreamStackBusOOB[34].pe__sys__thisSynchronized          ), 
        .pe34__sys__ready              ( DownstreamStackBusOOB[34].pe__sys__ready                     ), 
        .pe34__sys__complete           ( DownstreamStackBusOOB[34].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe35__allSynchronized    ( DownstreamStackBusOOB[35].cb_test.sys__pe__allSynchronized   ), 
        .pe35__sys__thisSynchronized   ( DownstreamStackBusOOB[35].pe__sys__thisSynchronized          ), 
        .pe35__sys__ready              ( DownstreamStackBusOOB[35].pe__sys__ready                     ), 
        .pe35__sys__complete           ( DownstreamStackBusOOB[35].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe36__allSynchronized    ( DownstreamStackBusOOB[36].cb_test.sys__pe__allSynchronized   ), 
        .pe36__sys__thisSynchronized   ( DownstreamStackBusOOB[36].pe__sys__thisSynchronized          ), 
        .pe36__sys__ready              ( DownstreamStackBusOOB[36].pe__sys__ready                     ), 
        .pe36__sys__complete           ( DownstreamStackBusOOB[36].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe37__allSynchronized    ( DownstreamStackBusOOB[37].cb_test.sys__pe__allSynchronized   ), 
        .pe37__sys__thisSynchronized   ( DownstreamStackBusOOB[37].pe__sys__thisSynchronized          ), 
        .pe37__sys__ready              ( DownstreamStackBusOOB[37].pe__sys__ready                     ), 
        .pe37__sys__complete           ( DownstreamStackBusOOB[37].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe38__allSynchronized    ( DownstreamStackBusOOB[38].cb_test.sys__pe__allSynchronized   ), 
        .pe38__sys__thisSynchronized   ( DownstreamStackBusOOB[38].pe__sys__thisSynchronized          ), 
        .pe38__sys__ready              ( DownstreamStackBusOOB[38].pe__sys__ready                     ), 
        .pe38__sys__complete           ( DownstreamStackBusOOB[38].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe39__allSynchronized    ( DownstreamStackBusOOB[39].cb_test.sys__pe__allSynchronized   ), 
        .pe39__sys__thisSynchronized   ( DownstreamStackBusOOB[39].pe__sys__thisSynchronized          ), 
        .pe39__sys__ready              ( DownstreamStackBusOOB[39].pe__sys__ready                     ), 
        .pe39__sys__complete           ( DownstreamStackBusOOB[39].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe40__allSynchronized    ( DownstreamStackBusOOB[40].cb_test.sys__pe__allSynchronized   ), 
        .pe40__sys__thisSynchronized   ( DownstreamStackBusOOB[40].pe__sys__thisSynchronized          ), 
        .pe40__sys__ready              ( DownstreamStackBusOOB[40].pe__sys__ready                     ), 
        .pe40__sys__complete           ( DownstreamStackBusOOB[40].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe41__allSynchronized    ( DownstreamStackBusOOB[41].cb_test.sys__pe__allSynchronized   ), 
        .pe41__sys__thisSynchronized   ( DownstreamStackBusOOB[41].pe__sys__thisSynchronized          ), 
        .pe41__sys__ready              ( DownstreamStackBusOOB[41].pe__sys__ready                     ), 
        .pe41__sys__complete           ( DownstreamStackBusOOB[41].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe42__allSynchronized    ( DownstreamStackBusOOB[42].cb_test.sys__pe__allSynchronized   ), 
        .pe42__sys__thisSynchronized   ( DownstreamStackBusOOB[42].pe__sys__thisSynchronized          ), 
        .pe42__sys__ready              ( DownstreamStackBusOOB[42].pe__sys__ready                     ), 
        .pe42__sys__complete           ( DownstreamStackBusOOB[42].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe43__allSynchronized    ( DownstreamStackBusOOB[43].cb_test.sys__pe__allSynchronized   ), 
        .pe43__sys__thisSynchronized   ( DownstreamStackBusOOB[43].pe__sys__thisSynchronized          ), 
        .pe43__sys__ready              ( DownstreamStackBusOOB[43].pe__sys__ready                     ), 
        .pe43__sys__complete           ( DownstreamStackBusOOB[43].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe44__allSynchronized    ( DownstreamStackBusOOB[44].cb_test.sys__pe__allSynchronized   ), 
        .pe44__sys__thisSynchronized   ( DownstreamStackBusOOB[44].pe__sys__thisSynchronized          ), 
        .pe44__sys__ready              ( DownstreamStackBusOOB[44].pe__sys__ready                     ), 
        .pe44__sys__complete           ( DownstreamStackBusOOB[44].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe45__allSynchronized    ( DownstreamStackBusOOB[45].cb_test.sys__pe__allSynchronized   ), 
        .pe45__sys__thisSynchronized   ( DownstreamStackBusOOB[45].pe__sys__thisSynchronized          ), 
        .pe45__sys__ready              ( DownstreamStackBusOOB[45].pe__sys__ready                     ), 
        .pe45__sys__complete           ( DownstreamStackBusOOB[45].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe46__allSynchronized    ( DownstreamStackBusOOB[46].cb_test.sys__pe__allSynchronized   ), 
        .pe46__sys__thisSynchronized   ( DownstreamStackBusOOB[46].pe__sys__thisSynchronized          ), 
        .pe46__sys__ready              ( DownstreamStackBusOOB[46].pe__sys__ready                     ), 
        .pe46__sys__complete           ( DownstreamStackBusOOB[46].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe47__allSynchronized    ( DownstreamStackBusOOB[47].cb_test.sys__pe__allSynchronized   ), 
        .pe47__sys__thisSynchronized   ( DownstreamStackBusOOB[47].pe__sys__thisSynchronized          ), 
        .pe47__sys__ready              ( DownstreamStackBusOOB[47].pe__sys__ready                     ), 
        .pe47__sys__complete           ( DownstreamStackBusOOB[47].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe48__allSynchronized    ( DownstreamStackBusOOB[48].cb_test.sys__pe__allSynchronized   ), 
        .pe48__sys__thisSynchronized   ( DownstreamStackBusOOB[48].pe__sys__thisSynchronized          ), 
        .pe48__sys__ready              ( DownstreamStackBusOOB[48].pe__sys__ready                     ), 
        .pe48__sys__complete           ( DownstreamStackBusOOB[48].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe49__allSynchronized    ( DownstreamStackBusOOB[49].cb_test.sys__pe__allSynchronized   ), 
        .pe49__sys__thisSynchronized   ( DownstreamStackBusOOB[49].pe__sys__thisSynchronized          ), 
        .pe49__sys__ready              ( DownstreamStackBusOOB[49].pe__sys__ready                     ), 
        .pe49__sys__complete           ( DownstreamStackBusOOB[49].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe50__allSynchronized    ( DownstreamStackBusOOB[50].cb_test.sys__pe__allSynchronized   ), 
        .pe50__sys__thisSynchronized   ( DownstreamStackBusOOB[50].pe__sys__thisSynchronized          ), 
        .pe50__sys__ready              ( DownstreamStackBusOOB[50].pe__sys__ready                     ), 
        .pe50__sys__complete           ( DownstreamStackBusOOB[50].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe51__allSynchronized    ( DownstreamStackBusOOB[51].cb_test.sys__pe__allSynchronized   ), 
        .pe51__sys__thisSynchronized   ( DownstreamStackBusOOB[51].pe__sys__thisSynchronized          ), 
        .pe51__sys__ready              ( DownstreamStackBusOOB[51].pe__sys__ready                     ), 
        .pe51__sys__complete           ( DownstreamStackBusOOB[51].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe52__allSynchronized    ( DownstreamStackBusOOB[52].cb_test.sys__pe__allSynchronized   ), 
        .pe52__sys__thisSynchronized   ( DownstreamStackBusOOB[52].pe__sys__thisSynchronized          ), 
        .pe52__sys__ready              ( DownstreamStackBusOOB[52].pe__sys__ready                     ), 
        .pe52__sys__complete           ( DownstreamStackBusOOB[52].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe53__allSynchronized    ( DownstreamStackBusOOB[53].cb_test.sys__pe__allSynchronized   ), 
        .pe53__sys__thisSynchronized   ( DownstreamStackBusOOB[53].pe__sys__thisSynchronized          ), 
        .pe53__sys__ready              ( DownstreamStackBusOOB[53].pe__sys__ready                     ), 
        .pe53__sys__complete           ( DownstreamStackBusOOB[53].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe54__allSynchronized    ( DownstreamStackBusOOB[54].cb_test.sys__pe__allSynchronized   ), 
        .pe54__sys__thisSynchronized   ( DownstreamStackBusOOB[54].pe__sys__thisSynchronized          ), 
        .pe54__sys__ready              ( DownstreamStackBusOOB[54].pe__sys__ready                     ), 
        .pe54__sys__complete           ( DownstreamStackBusOOB[54].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe55__allSynchronized    ( DownstreamStackBusOOB[55].cb_test.sys__pe__allSynchronized   ), 
        .pe55__sys__thisSynchronized   ( DownstreamStackBusOOB[55].pe__sys__thisSynchronized          ), 
        .pe55__sys__ready              ( DownstreamStackBusOOB[55].pe__sys__ready                     ), 
        .pe55__sys__complete           ( DownstreamStackBusOOB[55].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe56__allSynchronized    ( DownstreamStackBusOOB[56].cb_test.sys__pe__allSynchronized   ), 
        .pe56__sys__thisSynchronized   ( DownstreamStackBusOOB[56].pe__sys__thisSynchronized          ), 
        .pe56__sys__ready              ( DownstreamStackBusOOB[56].pe__sys__ready                     ), 
        .pe56__sys__complete           ( DownstreamStackBusOOB[56].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe57__allSynchronized    ( DownstreamStackBusOOB[57].cb_test.sys__pe__allSynchronized   ), 
        .pe57__sys__thisSynchronized   ( DownstreamStackBusOOB[57].pe__sys__thisSynchronized          ), 
        .pe57__sys__ready              ( DownstreamStackBusOOB[57].pe__sys__ready                     ), 
        .pe57__sys__complete           ( DownstreamStackBusOOB[57].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe58__allSynchronized    ( DownstreamStackBusOOB[58].cb_test.sys__pe__allSynchronized   ), 
        .pe58__sys__thisSynchronized   ( DownstreamStackBusOOB[58].pe__sys__thisSynchronized          ), 
        .pe58__sys__ready              ( DownstreamStackBusOOB[58].pe__sys__ready                     ), 
        .pe58__sys__complete           ( DownstreamStackBusOOB[58].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe59__allSynchronized    ( DownstreamStackBusOOB[59].cb_test.sys__pe__allSynchronized   ), 
        .pe59__sys__thisSynchronized   ( DownstreamStackBusOOB[59].pe__sys__thisSynchronized          ), 
        .pe59__sys__ready              ( DownstreamStackBusOOB[59].pe__sys__ready                     ), 
        .pe59__sys__complete           ( DownstreamStackBusOOB[59].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe60__allSynchronized    ( DownstreamStackBusOOB[60].cb_test.sys__pe__allSynchronized   ), 
        .pe60__sys__thisSynchronized   ( DownstreamStackBusOOB[60].pe__sys__thisSynchronized          ), 
        .pe60__sys__ready              ( DownstreamStackBusOOB[60].pe__sys__ready                     ), 
        .pe60__sys__complete           ( DownstreamStackBusOOB[60].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe61__allSynchronized    ( DownstreamStackBusOOB[61].cb_test.sys__pe__allSynchronized   ), 
        .pe61__sys__thisSynchronized   ( DownstreamStackBusOOB[61].pe__sys__thisSynchronized          ), 
        .pe61__sys__ready              ( DownstreamStackBusOOB[61].pe__sys__ready                     ), 
        .pe61__sys__complete           ( DownstreamStackBusOOB[61].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe62__allSynchronized    ( DownstreamStackBusOOB[62].cb_test.sys__pe__allSynchronized   ), 
        .pe62__sys__thisSynchronized   ( DownstreamStackBusOOB[62].pe__sys__thisSynchronized          ), 
        .pe62__sys__ready              ( DownstreamStackBusOOB[62].pe__sys__ready                     ), 
        .pe62__sys__complete           ( DownstreamStackBusOOB[62].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe63__allSynchronized    ( DownstreamStackBusOOB[63].cb_test.sys__pe__allSynchronized   ), 
        .pe63__sys__thisSynchronized   ( DownstreamStackBusOOB[63].pe__sys__thisSynchronized          ), 
        .pe63__sys__ready              ( DownstreamStackBusOOB[63].pe__sys__ready                     ), 
        .pe63__sys__complete           ( DownstreamStackBusOOB[63].pe__sys__complete                  ), 
