`ifndef _simd_core_vh
`define _simd_core_vh

/*****************************************************************

    File name   : simd_core.vh
    Author      : Lee Baker
    Affiliation : North Carolina State University, Raleigh, NC
    Date        : June 2017
    email       : lbbaker@ncsu.edu

*****************************************************************/





//------------------------------------------------------------------------------------------------------------



`endif
