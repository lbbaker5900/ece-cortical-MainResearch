
  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[0].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[0].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[0].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[0].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[0].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[0].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[0].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[0].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[1].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[1].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[1].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[1].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[1].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[1].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[1].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[1].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[2].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[2].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[2].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[2].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[2].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[2].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[2].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[2].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[3].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[3].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[3].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[3].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[3].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[3].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[3].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[3].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[4].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[4].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[4].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[4].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[4].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[4].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[4].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[4].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[5].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[5].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[5].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[5].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[5].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[5].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[5].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[5].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[6].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[6].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[6].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[6].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[6].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[6].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[6].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[6].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[7].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[7].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[7].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[7].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[7].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[7].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[7].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[7].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[8].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[8].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[8].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[8].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[8].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[8].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[8].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[8].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[9].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[9].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[9].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[9].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[9].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[9].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[9].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[9].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[10].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[10].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[10].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[10].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[10].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[10].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[10].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[10].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[11].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[11].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[11].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[11].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[11].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[11].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[11].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[11].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[12].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[12].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[12].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[12].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[12].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[12].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[12].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[12].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[13].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[13].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[13].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[13].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[13].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[13].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[13].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[13].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[14].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[14].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[14].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[14].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[14].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[14].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[14].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[14].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[15].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[15].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[15].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[15].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[15].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[15].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[15].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[15].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[16].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[16].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[16].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[16].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[16].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[16].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[16].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[16].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[17].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[17].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[17].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[17].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[17].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[17].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[17].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[17].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[18].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[18].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[18].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[18].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[18].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[18].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[18].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[18].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[19].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[19].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[19].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[19].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[19].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[19].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[19].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[19].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[20].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[20].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[20].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[20].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[20].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[20].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[20].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[20].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[21].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[21].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[21].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[21].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[21].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[21].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[21].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[21].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[22].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[22].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[22].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[22].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[22].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[22].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[22].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[22].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[23].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[23].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[23].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[23].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[23].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[23].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[23].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[23].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[24].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[24].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[24].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[24].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[24].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[24].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[24].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[24].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[25].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[25].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[25].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[25].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[25].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[25].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[25].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[25].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[26].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[26].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[26].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[26].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[26].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[26].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[26].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[26].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[27].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[27].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[27].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[27].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[27].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[27].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[27].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[27].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[28].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[28].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[28].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[28].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[28].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[28].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[28].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[28].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[29].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[29].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[29].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[29].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[29].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[29].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[29].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[29].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[30].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[30].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[30].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[30].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[30].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[30].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[30].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[30].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[31].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[31].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[31].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[31].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[31].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[31].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[31].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[31].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[32].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[32].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[32].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[32].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[32].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[32].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[32].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[32].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[33].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[33].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[33].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[33].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[33].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[33].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[33].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[33].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[34].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[34].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[34].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[34].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[34].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[34].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[34].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[34].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[35].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[35].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[35].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[35].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[35].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[35].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[35].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[35].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[36].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[36].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[36].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[36].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[36].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[36].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[36].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[36].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[37].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[37].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[37].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[37].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[37].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[37].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[37].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[37].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[38].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[38].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[38].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[38].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[38].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[38].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[38].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[38].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[39].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[39].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[39].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[39].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[39].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[39].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[39].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[39].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[40].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[40].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[40].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[40].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[40].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[40].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[40].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[40].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[41].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[41].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[41].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[41].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[41].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[41].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[41].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[41].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[42].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[42].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[42].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[42].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[42].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[42].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[42].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[42].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[43].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[43].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[43].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[43].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[43].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[43].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[43].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[43].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[44].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[44].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[44].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[44].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[44].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[44].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[44].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[44].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[45].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[45].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[45].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[45].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[45].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[45].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[45].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[45].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[46].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[46].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[46].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[46].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[46].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[46].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[46].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[46].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[47].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[47].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[47].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[47].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[47].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[47].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[47].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[47].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[48].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[48].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[48].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[48].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[48].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[48].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[48].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[48].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[49].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[49].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[49].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[49].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[49].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[49].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[49].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[49].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[50].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[50].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[50].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[50].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[50].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[50].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[50].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[50].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[51].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[51].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[51].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[51].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[51].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[51].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[51].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[51].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[52].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[52].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[52].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[52].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[52].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[52].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[52].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[52].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[53].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[53].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[53].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[53].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[53].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[53].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[53].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[53].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[54].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[54].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[54].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[54].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[54].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[54].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[54].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[54].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[55].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[55].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[55].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[55].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[55].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[55].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[55].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[55].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[56].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[56].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[56].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[56].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[56].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[56].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[56].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[56].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[57].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[57].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[57].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[57].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[57].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[57].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[57].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[57].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[58].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[58].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[58].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[58].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[58].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[58].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[58].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[58].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[59].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[59].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[59].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[59].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[59].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[59].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[59].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[59].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[60].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[60].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[60].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[60].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[60].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[60].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[60].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[60].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[61].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[61].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[61].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[61].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[61].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[61].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[61].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[61].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[62].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[62].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[62].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[62].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[62].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[62].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[62].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[62].sys__mgr__complete           ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[63].mgr__sys__allSynchronized   =   DownstreamStackBusOOB[63].sys__pe__allSynchronized                      ; 
  assign DownstreamStackBusOOB[63].pe__sys__thisSynchronized                     =  system_inst.manager_array_inst.mgr_inst[63].sys__mgr__thisSynchronized   ; 
  assign DownstreamStackBusOOB[63].pe__sys__ready                                =  system_inst.manager_array_inst.mgr_inst[63].sys__mgr__ready              ; 
  assign DownstreamStackBusOOB[63].pe__sys__complete                             =  system_inst.manager_array_inst.mgr_inst[63].sys__mgr__complete           ; 
