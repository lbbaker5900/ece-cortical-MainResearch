
  assign   pe_inst[0].sys__pe__allSynchronized    =  sys__pe0__allSynchronized                ;
  assign   pe0__sys__thisSynchronized             =  pe_inst[0].pe__sys__thisSynchronized     ;
  assign   pe0__sys__ready                        =  pe_inst[0].pe__sys__ready                ;
  assign   pe0__sys__complete                     =  pe_inst[0].pe__sys__complete             ;
  assign   pe_inst[0].std__pe__oob_cntl           =  std__pe0__oob_cntl                       ;
  assign   pe_inst[0].std__pe__oob_valid          =  std__pe0__oob_valid                      ;
  assign   pe0__std__oob_ready                    =  pe_inst[0].pe__std__oob_ready            ;
  assign   pe_inst[0].std__pe__oob_type           =  std__pe0__oob_type                       ;
  assign   pe_inst[0].std__pe__oob_data           =  std__pe0__oob_data                       ;
  assign   pe_inst[1].sys__pe__allSynchronized    =  sys__pe1__allSynchronized                ;
  assign   pe1__sys__thisSynchronized             =  pe_inst[1].pe__sys__thisSynchronized     ;
  assign   pe1__sys__ready                        =  pe_inst[1].pe__sys__ready                ;
  assign   pe1__sys__complete                     =  pe_inst[1].pe__sys__complete             ;
  assign   pe_inst[1].std__pe__oob_cntl           =  std__pe1__oob_cntl                       ;
  assign   pe_inst[1].std__pe__oob_valid          =  std__pe1__oob_valid                      ;
  assign   pe1__std__oob_ready                    =  pe_inst[1].pe__std__oob_ready            ;
  assign   pe_inst[1].std__pe__oob_type           =  std__pe1__oob_type                       ;
  assign   pe_inst[1].std__pe__oob_data           =  std__pe1__oob_data                       ;
  assign   pe_inst[2].sys__pe__allSynchronized    =  sys__pe2__allSynchronized                ;
  assign   pe2__sys__thisSynchronized             =  pe_inst[2].pe__sys__thisSynchronized     ;
  assign   pe2__sys__ready                        =  pe_inst[2].pe__sys__ready                ;
  assign   pe2__sys__complete                     =  pe_inst[2].pe__sys__complete             ;
  assign   pe_inst[2].std__pe__oob_cntl           =  std__pe2__oob_cntl                       ;
  assign   pe_inst[2].std__pe__oob_valid          =  std__pe2__oob_valid                      ;
  assign   pe2__std__oob_ready                    =  pe_inst[2].pe__std__oob_ready            ;
  assign   pe_inst[2].std__pe__oob_type           =  std__pe2__oob_type                       ;
  assign   pe_inst[2].std__pe__oob_data           =  std__pe2__oob_data                       ;
  assign   pe_inst[3].sys__pe__allSynchronized    =  sys__pe3__allSynchronized                ;
  assign   pe3__sys__thisSynchronized             =  pe_inst[3].pe__sys__thisSynchronized     ;
  assign   pe3__sys__ready                        =  pe_inst[3].pe__sys__ready                ;
  assign   pe3__sys__complete                     =  pe_inst[3].pe__sys__complete             ;
  assign   pe_inst[3].std__pe__oob_cntl           =  std__pe3__oob_cntl                       ;
  assign   pe_inst[3].std__pe__oob_valid          =  std__pe3__oob_valid                      ;
  assign   pe3__std__oob_ready                    =  pe_inst[3].pe__std__oob_ready            ;
  assign   pe_inst[3].std__pe__oob_type           =  std__pe3__oob_type                       ;
  assign   pe_inst[3].std__pe__oob_data           =  std__pe3__oob_data                       ;
