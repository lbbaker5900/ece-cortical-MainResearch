
  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe0__peId                ;
  input                                         sys__pe0__allSynchronized     ;
  output                                        pe0__sys__thisSynchronized    ;
  output                                        pe0__sys__ready               ;
  output                                        pe0__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe0__oob_cntl            ;
  input                                         std__pe0__oob_valid           ;
  output                                        pe0__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe0__oob_type            ;
  output                                          pe0__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane0_strm0_data_mask   ;
  input                                           std__pe0__lane0_strm0_data_valid  ;

  output                                          pe0__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane0_strm1_data_mask   ;
  input                                           std__pe0__lane0_strm1_data_valid  ;

  output                                          pe0__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane1_strm0_data_mask   ;
  input                                           std__pe0__lane1_strm0_data_valid  ;

  output                                          pe0__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane1_strm1_data_mask   ;
  input                                           std__pe0__lane1_strm1_data_valid  ;

  output                                          pe0__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane2_strm0_data_mask   ;
  input                                           std__pe0__lane2_strm0_data_valid  ;

  output                                          pe0__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane2_strm1_data_mask   ;
  input                                           std__pe0__lane2_strm1_data_valid  ;

  output                                          pe0__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane3_strm0_data_mask   ;
  input                                           std__pe0__lane3_strm0_data_valid  ;

  output                                          pe0__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane3_strm1_data_mask   ;
  input                                           std__pe0__lane3_strm1_data_valid  ;

  output                                          pe0__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane4_strm0_data_mask   ;
  input                                           std__pe0__lane4_strm0_data_valid  ;

  output                                          pe0__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane4_strm1_data_mask   ;
  input                                           std__pe0__lane4_strm1_data_valid  ;

  output                                          pe0__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane5_strm0_data_mask   ;
  input                                           std__pe0__lane5_strm0_data_valid  ;

  output                                          pe0__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane5_strm1_data_mask   ;
  input                                           std__pe0__lane5_strm1_data_valid  ;

  output                                          pe0__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane6_strm0_data_mask   ;
  input                                           std__pe0__lane6_strm0_data_valid  ;

  output                                          pe0__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane6_strm1_data_mask   ;
  input                                           std__pe0__lane6_strm1_data_valid  ;

  output                                          pe0__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane7_strm0_data_mask   ;
  input                                           std__pe0__lane7_strm0_data_valid  ;

  output                                          pe0__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane7_strm1_data_mask   ;
  input                                           std__pe0__lane7_strm1_data_valid  ;

  output                                          pe0__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane8_strm0_data_mask   ;
  input                                           std__pe0__lane8_strm0_data_valid  ;

  output                                          pe0__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane8_strm1_data_mask   ;
  input                                           std__pe0__lane8_strm1_data_valid  ;

  output                                          pe0__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane9_strm0_data_mask   ;
  input                                           std__pe0__lane9_strm0_data_valid  ;

  output                                          pe0__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane9_strm1_data_mask   ;
  input                                           std__pe0__lane9_strm1_data_valid  ;

  output                                          pe0__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane10_strm0_data_mask   ;
  input                                           std__pe0__lane10_strm0_data_valid  ;

  output                                          pe0__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane10_strm1_data_mask   ;
  input                                           std__pe0__lane10_strm1_data_valid  ;

  output                                          pe0__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane11_strm0_data_mask   ;
  input                                           std__pe0__lane11_strm0_data_valid  ;

  output                                          pe0__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane11_strm1_data_mask   ;
  input                                           std__pe0__lane11_strm1_data_valid  ;

  output                                          pe0__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane12_strm0_data_mask   ;
  input                                           std__pe0__lane12_strm0_data_valid  ;

  output                                          pe0__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane12_strm1_data_mask   ;
  input                                           std__pe0__lane12_strm1_data_valid  ;

  output                                          pe0__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane13_strm0_data_mask   ;
  input                                           std__pe0__lane13_strm0_data_valid  ;

  output                                          pe0__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane13_strm1_data_mask   ;
  input                                           std__pe0__lane13_strm1_data_valid  ;

  output                                          pe0__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane14_strm0_data_mask   ;
  input                                           std__pe0__lane14_strm0_data_valid  ;

  output                                          pe0__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane14_strm1_data_mask   ;
  input                                           std__pe0__lane14_strm1_data_valid  ;

  output                                          pe0__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane15_strm0_data_mask   ;
  input                                           std__pe0__lane15_strm0_data_valid  ;

  output                                          pe0__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane15_strm1_data_mask   ;
  input                                           std__pe0__lane15_strm1_data_valid  ;

  output                                          pe0__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane16_strm0_data_mask   ;
  input                                           std__pe0__lane16_strm0_data_valid  ;

  output                                          pe0__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane16_strm1_data_mask   ;
  input                                           std__pe0__lane16_strm1_data_valid  ;

  output                                          pe0__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane17_strm0_data_mask   ;
  input                                           std__pe0__lane17_strm0_data_valid  ;

  output                                          pe0__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane17_strm1_data_mask   ;
  input                                           std__pe0__lane17_strm1_data_valid  ;

  output                                          pe0__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane18_strm0_data_mask   ;
  input                                           std__pe0__lane18_strm0_data_valid  ;

  output                                          pe0__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane18_strm1_data_mask   ;
  input                                           std__pe0__lane18_strm1_data_valid  ;

  output                                          pe0__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane19_strm0_data_mask   ;
  input                                           std__pe0__lane19_strm0_data_valid  ;

  output                                          pe0__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane19_strm1_data_mask   ;
  input                                           std__pe0__lane19_strm1_data_valid  ;

  output                                          pe0__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane20_strm0_data_mask   ;
  input                                           std__pe0__lane20_strm0_data_valid  ;

  output                                          pe0__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane20_strm1_data_mask   ;
  input                                           std__pe0__lane20_strm1_data_valid  ;

  output                                          pe0__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane21_strm0_data_mask   ;
  input                                           std__pe0__lane21_strm0_data_valid  ;

  output                                          pe0__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane21_strm1_data_mask   ;
  input                                           std__pe0__lane21_strm1_data_valid  ;

  output                                          pe0__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane22_strm0_data_mask   ;
  input                                           std__pe0__lane22_strm0_data_valid  ;

  output                                          pe0__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane22_strm1_data_mask   ;
  input                                           std__pe0__lane22_strm1_data_valid  ;

  output                                          pe0__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane23_strm0_data_mask   ;
  input                                           std__pe0__lane23_strm0_data_valid  ;

  output                                          pe0__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane23_strm1_data_mask   ;
  input                                           std__pe0__lane23_strm1_data_valid  ;

  output                                          pe0__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane24_strm0_data_mask   ;
  input                                           std__pe0__lane24_strm0_data_valid  ;

  output                                          pe0__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane24_strm1_data_mask   ;
  input                                           std__pe0__lane24_strm1_data_valid  ;

  output                                          pe0__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane25_strm0_data_mask   ;
  input                                           std__pe0__lane25_strm0_data_valid  ;

  output                                          pe0__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane25_strm1_data_mask   ;
  input                                           std__pe0__lane25_strm1_data_valid  ;

  output                                          pe0__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane26_strm0_data_mask   ;
  input                                           std__pe0__lane26_strm0_data_valid  ;

  output                                          pe0__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane26_strm1_data_mask   ;
  input                                           std__pe0__lane26_strm1_data_valid  ;

  output                                          pe0__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane27_strm0_data_mask   ;
  input                                           std__pe0__lane27_strm0_data_valid  ;

  output                                          pe0__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane27_strm1_data_mask   ;
  input                                           std__pe0__lane27_strm1_data_valid  ;

  output                                          pe0__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane28_strm0_data_mask   ;
  input                                           std__pe0__lane28_strm0_data_valid  ;

  output                                          pe0__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane28_strm1_data_mask   ;
  input                                           std__pe0__lane28_strm1_data_valid  ;

  output                                          pe0__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane29_strm0_data_mask   ;
  input                                           std__pe0__lane29_strm0_data_valid  ;

  output                                          pe0__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane29_strm1_data_mask   ;
  input                                           std__pe0__lane29_strm1_data_valid  ;

  output                                          pe0__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane30_strm0_data_mask   ;
  input                                           std__pe0__lane30_strm0_data_valid  ;

  output                                          pe0__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane30_strm1_data_mask   ;
  input                                           std__pe0__lane30_strm1_data_valid  ;

  output                                          pe0__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane31_strm0_data_mask   ;
  input                                           std__pe0__lane31_strm0_data_valid  ;

  output                                          pe0__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe0__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe0__lane31_strm1_data_mask   ;
  input                                           std__pe0__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe1__peId                ;
  input                                         sys__pe1__allSynchronized     ;
  output                                        pe1__sys__thisSynchronized    ;
  output                                        pe1__sys__ready               ;
  output                                        pe1__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe1__oob_cntl            ;
  input                                         std__pe1__oob_valid           ;
  output                                        pe1__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe1__oob_type            ;
  output                                          pe1__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane0_strm0_data_mask   ;
  input                                           std__pe1__lane0_strm0_data_valid  ;

  output                                          pe1__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane0_strm1_data_mask   ;
  input                                           std__pe1__lane0_strm1_data_valid  ;

  output                                          pe1__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane1_strm0_data_mask   ;
  input                                           std__pe1__lane1_strm0_data_valid  ;

  output                                          pe1__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane1_strm1_data_mask   ;
  input                                           std__pe1__lane1_strm1_data_valid  ;

  output                                          pe1__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane2_strm0_data_mask   ;
  input                                           std__pe1__lane2_strm0_data_valid  ;

  output                                          pe1__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane2_strm1_data_mask   ;
  input                                           std__pe1__lane2_strm1_data_valid  ;

  output                                          pe1__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane3_strm0_data_mask   ;
  input                                           std__pe1__lane3_strm0_data_valid  ;

  output                                          pe1__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane3_strm1_data_mask   ;
  input                                           std__pe1__lane3_strm1_data_valid  ;

  output                                          pe1__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane4_strm0_data_mask   ;
  input                                           std__pe1__lane4_strm0_data_valid  ;

  output                                          pe1__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane4_strm1_data_mask   ;
  input                                           std__pe1__lane4_strm1_data_valid  ;

  output                                          pe1__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane5_strm0_data_mask   ;
  input                                           std__pe1__lane5_strm0_data_valid  ;

  output                                          pe1__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane5_strm1_data_mask   ;
  input                                           std__pe1__lane5_strm1_data_valid  ;

  output                                          pe1__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane6_strm0_data_mask   ;
  input                                           std__pe1__lane6_strm0_data_valid  ;

  output                                          pe1__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane6_strm1_data_mask   ;
  input                                           std__pe1__lane6_strm1_data_valid  ;

  output                                          pe1__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane7_strm0_data_mask   ;
  input                                           std__pe1__lane7_strm0_data_valid  ;

  output                                          pe1__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane7_strm1_data_mask   ;
  input                                           std__pe1__lane7_strm1_data_valid  ;

  output                                          pe1__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane8_strm0_data_mask   ;
  input                                           std__pe1__lane8_strm0_data_valid  ;

  output                                          pe1__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane8_strm1_data_mask   ;
  input                                           std__pe1__lane8_strm1_data_valid  ;

  output                                          pe1__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane9_strm0_data_mask   ;
  input                                           std__pe1__lane9_strm0_data_valid  ;

  output                                          pe1__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane9_strm1_data_mask   ;
  input                                           std__pe1__lane9_strm1_data_valid  ;

  output                                          pe1__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane10_strm0_data_mask   ;
  input                                           std__pe1__lane10_strm0_data_valid  ;

  output                                          pe1__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane10_strm1_data_mask   ;
  input                                           std__pe1__lane10_strm1_data_valid  ;

  output                                          pe1__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane11_strm0_data_mask   ;
  input                                           std__pe1__lane11_strm0_data_valid  ;

  output                                          pe1__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane11_strm1_data_mask   ;
  input                                           std__pe1__lane11_strm1_data_valid  ;

  output                                          pe1__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane12_strm0_data_mask   ;
  input                                           std__pe1__lane12_strm0_data_valid  ;

  output                                          pe1__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane12_strm1_data_mask   ;
  input                                           std__pe1__lane12_strm1_data_valid  ;

  output                                          pe1__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane13_strm0_data_mask   ;
  input                                           std__pe1__lane13_strm0_data_valid  ;

  output                                          pe1__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane13_strm1_data_mask   ;
  input                                           std__pe1__lane13_strm1_data_valid  ;

  output                                          pe1__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane14_strm0_data_mask   ;
  input                                           std__pe1__lane14_strm0_data_valid  ;

  output                                          pe1__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane14_strm1_data_mask   ;
  input                                           std__pe1__lane14_strm1_data_valid  ;

  output                                          pe1__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane15_strm0_data_mask   ;
  input                                           std__pe1__lane15_strm0_data_valid  ;

  output                                          pe1__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane15_strm1_data_mask   ;
  input                                           std__pe1__lane15_strm1_data_valid  ;

  output                                          pe1__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane16_strm0_data_mask   ;
  input                                           std__pe1__lane16_strm0_data_valid  ;

  output                                          pe1__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane16_strm1_data_mask   ;
  input                                           std__pe1__lane16_strm1_data_valid  ;

  output                                          pe1__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane17_strm0_data_mask   ;
  input                                           std__pe1__lane17_strm0_data_valid  ;

  output                                          pe1__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane17_strm1_data_mask   ;
  input                                           std__pe1__lane17_strm1_data_valid  ;

  output                                          pe1__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane18_strm0_data_mask   ;
  input                                           std__pe1__lane18_strm0_data_valid  ;

  output                                          pe1__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane18_strm1_data_mask   ;
  input                                           std__pe1__lane18_strm1_data_valid  ;

  output                                          pe1__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane19_strm0_data_mask   ;
  input                                           std__pe1__lane19_strm0_data_valid  ;

  output                                          pe1__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane19_strm1_data_mask   ;
  input                                           std__pe1__lane19_strm1_data_valid  ;

  output                                          pe1__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane20_strm0_data_mask   ;
  input                                           std__pe1__lane20_strm0_data_valid  ;

  output                                          pe1__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane20_strm1_data_mask   ;
  input                                           std__pe1__lane20_strm1_data_valid  ;

  output                                          pe1__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane21_strm0_data_mask   ;
  input                                           std__pe1__lane21_strm0_data_valid  ;

  output                                          pe1__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane21_strm1_data_mask   ;
  input                                           std__pe1__lane21_strm1_data_valid  ;

  output                                          pe1__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane22_strm0_data_mask   ;
  input                                           std__pe1__lane22_strm0_data_valid  ;

  output                                          pe1__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane22_strm1_data_mask   ;
  input                                           std__pe1__lane22_strm1_data_valid  ;

  output                                          pe1__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane23_strm0_data_mask   ;
  input                                           std__pe1__lane23_strm0_data_valid  ;

  output                                          pe1__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane23_strm1_data_mask   ;
  input                                           std__pe1__lane23_strm1_data_valid  ;

  output                                          pe1__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane24_strm0_data_mask   ;
  input                                           std__pe1__lane24_strm0_data_valid  ;

  output                                          pe1__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane24_strm1_data_mask   ;
  input                                           std__pe1__lane24_strm1_data_valid  ;

  output                                          pe1__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane25_strm0_data_mask   ;
  input                                           std__pe1__lane25_strm0_data_valid  ;

  output                                          pe1__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane25_strm1_data_mask   ;
  input                                           std__pe1__lane25_strm1_data_valid  ;

  output                                          pe1__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane26_strm0_data_mask   ;
  input                                           std__pe1__lane26_strm0_data_valid  ;

  output                                          pe1__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane26_strm1_data_mask   ;
  input                                           std__pe1__lane26_strm1_data_valid  ;

  output                                          pe1__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane27_strm0_data_mask   ;
  input                                           std__pe1__lane27_strm0_data_valid  ;

  output                                          pe1__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane27_strm1_data_mask   ;
  input                                           std__pe1__lane27_strm1_data_valid  ;

  output                                          pe1__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane28_strm0_data_mask   ;
  input                                           std__pe1__lane28_strm0_data_valid  ;

  output                                          pe1__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane28_strm1_data_mask   ;
  input                                           std__pe1__lane28_strm1_data_valid  ;

  output                                          pe1__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane29_strm0_data_mask   ;
  input                                           std__pe1__lane29_strm0_data_valid  ;

  output                                          pe1__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane29_strm1_data_mask   ;
  input                                           std__pe1__lane29_strm1_data_valid  ;

  output                                          pe1__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane30_strm0_data_mask   ;
  input                                           std__pe1__lane30_strm0_data_valid  ;

  output                                          pe1__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane30_strm1_data_mask   ;
  input                                           std__pe1__lane30_strm1_data_valid  ;

  output                                          pe1__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane31_strm0_data_mask   ;
  input                                           std__pe1__lane31_strm0_data_valid  ;

  output                                          pe1__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe1__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe1__lane31_strm1_data_mask   ;
  input                                           std__pe1__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe2__peId                ;
  input                                         sys__pe2__allSynchronized     ;
  output                                        pe2__sys__thisSynchronized    ;
  output                                        pe2__sys__ready               ;
  output                                        pe2__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe2__oob_cntl            ;
  input                                         std__pe2__oob_valid           ;
  output                                        pe2__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe2__oob_type            ;
  output                                          pe2__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane0_strm0_data_mask   ;
  input                                           std__pe2__lane0_strm0_data_valid  ;

  output                                          pe2__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane0_strm1_data_mask   ;
  input                                           std__pe2__lane0_strm1_data_valid  ;

  output                                          pe2__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane1_strm0_data_mask   ;
  input                                           std__pe2__lane1_strm0_data_valid  ;

  output                                          pe2__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane1_strm1_data_mask   ;
  input                                           std__pe2__lane1_strm1_data_valid  ;

  output                                          pe2__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane2_strm0_data_mask   ;
  input                                           std__pe2__lane2_strm0_data_valid  ;

  output                                          pe2__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane2_strm1_data_mask   ;
  input                                           std__pe2__lane2_strm1_data_valid  ;

  output                                          pe2__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane3_strm0_data_mask   ;
  input                                           std__pe2__lane3_strm0_data_valid  ;

  output                                          pe2__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane3_strm1_data_mask   ;
  input                                           std__pe2__lane3_strm1_data_valid  ;

  output                                          pe2__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane4_strm0_data_mask   ;
  input                                           std__pe2__lane4_strm0_data_valid  ;

  output                                          pe2__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane4_strm1_data_mask   ;
  input                                           std__pe2__lane4_strm1_data_valid  ;

  output                                          pe2__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane5_strm0_data_mask   ;
  input                                           std__pe2__lane5_strm0_data_valid  ;

  output                                          pe2__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane5_strm1_data_mask   ;
  input                                           std__pe2__lane5_strm1_data_valid  ;

  output                                          pe2__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane6_strm0_data_mask   ;
  input                                           std__pe2__lane6_strm0_data_valid  ;

  output                                          pe2__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane6_strm1_data_mask   ;
  input                                           std__pe2__lane6_strm1_data_valid  ;

  output                                          pe2__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane7_strm0_data_mask   ;
  input                                           std__pe2__lane7_strm0_data_valid  ;

  output                                          pe2__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane7_strm1_data_mask   ;
  input                                           std__pe2__lane7_strm1_data_valid  ;

  output                                          pe2__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane8_strm0_data_mask   ;
  input                                           std__pe2__lane8_strm0_data_valid  ;

  output                                          pe2__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane8_strm1_data_mask   ;
  input                                           std__pe2__lane8_strm1_data_valid  ;

  output                                          pe2__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane9_strm0_data_mask   ;
  input                                           std__pe2__lane9_strm0_data_valid  ;

  output                                          pe2__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane9_strm1_data_mask   ;
  input                                           std__pe2__lane9_strm1_data_valid  ;

  output                                          pe2__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane10_strm0_data_mask   ;
  input                                           std__pe2__lane10_strm0_data_valid  ;

  output                                          pe2__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane10_strm1_data_mask   ;
  input                                           std__pe2__lane10_strm1_data_valid  ;

  output                                          pe2__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane11_strm0_data_mask   ;
  input                                           std__pe2__lane11_strm0_data_valid  ;

  output                                          pe2__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane11_strm1_data_mask   ;
  input                                           std__pe2__lane11_strm1_data_valid  ;

  output                                          pe2__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane12_strm0_data_mask   ;
  input                                           std__pe2__lane12_strm0_data_valid  ;

  output                                          pe2__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane12_strm1_data_mask   ;
  input                                           std__pe2__lane12_strm1_data_valid  ;

  output                                          pe2__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane13_strm0_data_mask   ;
  input                                           std__pe2__lane13_strm0_data_valid  ;

  output                                          pe2__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane13_strm1_data_mask   ;
  input                                           std__pe2__lane13_strm1_data_valid  ;

  output                                          pe2__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane14_strm0_data_mask   ;
  input                                           std__pe2__lane14_strm0_data_valid  ;

  output                                          pe2__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane14_strm1_data_mask   ;
  input                                           std__pe2__lane14_strm1_data_valid  ;

  output                                          pe2__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane15_strm0_data_mask   ;
  input                                           std__pe2__lane15_strm0_data_valid  ;

  output                                          pe2__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane15_strm1_data_mask   ;
  input                                           std__pe2__lane15_strm1_data_valid  ;

  output                                          pe2__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane16_strm0_data_mask   ;
  input                                           std__pe2__lane16_strm0_data_valid  ;

  output                                          pe2__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane16_strm1_data_mask   ;
  input                                           std__pe2__lane16_strm1_data_valid  ;

  output                                          pe2__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane17_strm0_data_mask   ;
  input                                           std__pe2__lane17_strm0_data_valid  ;

  output                                          pe2__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane17_strm1_data_mask   ;
  input                                           std__pe2__lane17_strm1_data_valid  ;

  output                                          pe2__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane18_strm0_data_mask   ;
  input                                           std__pe2__lane18_strm0_data_valid  ;

  output                                          pe2__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane18_strm1_data_mask   ;
  input                                           std__pe2__lane18_strm1_data_valid  ;

  output                                          pe2__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane19_strm0_data_mask   ;
  input                                           std__pe2__lane19_strm0_data_valid  ;

  output                                          pe2__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane19_strm1_data_mask   ;
  input                                           std__pe2__lane19_strm1_data_valid  ;

  output                                          pe2__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane20_strm0_data_mask   ;
  input                                           std__pe2__lane20_strm0_data_valid  ;

  output                                          pe2__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane20_strm1_data_mask   ;
  input                                           std__pe2__lane20_strm1_data_valid  ;

  output                                          pe2__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane21_strm0_data_mask   ;
  input                                           std__pe2__lane21_strm0_data_valid  ;

  output                                          pe2__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane21_strm1_data_mask   ;
  input                                           std__pe2__lane21_strm1_data_valid  ;

  output                                          pe2__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane22_strm0_data_mask   ;
  input                                           std__pe2__lane22_strm0_data_valid  ;

  output                                          pe2__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane22_strm1_data_mask   ;
  input                                           std__pe2__lane22_strm1_data_valid  ;

  output                                          pe2__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane23_strm0_data_mask   ;
  input                                           std__pe2__lane23_strm0_data_valid  ;

  output                                          pe2__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane23_strm1_data_mask   ;
  input                                           std__pe2__lane23_strm1_data_valid  ;

  output                                          pe2__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane24_strm0_data_mask   ;
  input                                           std__pe2__lane24_strm0_data_valid  ;

  output                                          pe2__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane24_strm1_data_mask   ;
  input                                           std__pe2__lane24_strm1_data_valid  ;

  output                                          pe2__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane25_strm0_data_mask   ;
  input                                           std__pe2__lane25_strm0_data_valid  ;

  output                                          pe2__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane25_strm1_data_mask   ;
  input                                           std__pe2__lane25_strm1_data_valid  ;

  output                                          pe2__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane26_strm0_data_mask   ;
  input                                           std__pe2__lane26_strm0_data_valid  ;

  output                                          pe2__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane26_strm1_data_mask   ;
  input                                           std__pe2__lane26_strm1_data_valid  ;

  output                                          pe2__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane27_strm0_data_mask   ;
  input                                           std__pe2__lane27_strm0_data_valid  ;

  output                                          pe2__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane27_strm1_data_mask   ;
  input                                           std__pe2__lane27_strm1_data_valid  ;

  output                                          pe2__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane28_strm0_data_mask   ;
  input                                           std__pe2__lane28_strm0_data_valid  ;

  output                                          pe2__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane28_strm1_data_mask   ;
  input                                           std__pe2__lane28_strm1_data_valid  ;

  output                                          pe2__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane29_strm0_data_mask   ;
  input                                           std__pe2__lane29_strm0_data_valid  ;

  output                                          pe2__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane29_strm1_data_mask   ;
  input                                           std__pe2__lane29_strm1_data_valid  ;

  output                                          pe2__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane30_strm0_data_mask   ;
  input                                           std__pe2__lane30_strm0_data_valid  ;

  output                                          pe2__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane30_strm1_data_mask   ;
  input                                           std__pe2__lane30_strm1_data_valid  ;

  output                                          pe2__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane31_strm0_data_mask   ;
  input                                           std__pe2__lane31_strm0_data_valid  ;

  output                                          pe2__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe2__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe2__lane31_strm1_data_mask   ;
  input                                           std__pe2__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe3__peId                ;
  input                                         sys__pe3__allSynchronized     ;
  output                                        pe3__sys__thisSynchronized    ;
  output                                        pe3__sys__ready               ;
  output                                        pe3__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe3__oob_cntl            ;
  input                                         std__pe3__oob_valid           ;
  output                                        pe3__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe3__oob_type            ;
  output                                          pe3__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane0_strm0_data_mask   ;
  input                                           std__pe3__lane0_strm0_data_valid  ;

  output                                          pe3__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane0_strm1_data_mask   ;
  input                                           std__pe3__lane0_strm1_data_valid  ;

  output                                          pe3__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane1_strm0_data_mask   ;
  input                                           std__pe3__lane1_strm0_data_valid  ;

  output                                          pe3__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane1_strm1_data_mask   ;
  input                                           std__pe3__lane1_strm1_data_valid  ;

  output                                          pe3__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane2_strm0_data_mask   ;
  input                                           std__pe3__lane2_strm0_data_valid  ;

  output                                          pe3__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane2_strm1_data_mask   ;
  input                                           std__pe3__lane2_strm1_data_valid  ;

  output                                          pe3__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane3_strm0_data_mask   ;
  input                                           std__pe3__lane3_strm0_data_valid  ;

  output                                          pe3__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane3_strm1_data_mask   ;
  input                                           std__pe3__lane3_strm1_data_valid  ;

  output                                          pe3__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane4_strm0_data_mask   ;
  input                                           std__pe3__lane4_strm0_data_valid  ;

  output                                          pe3__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane4_strm1_data_mask   ;
  input                                           std__pe3__lane4_strm1_data_valid  ;

  output                                          pe3__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane5_strm0_data_mask   ;
  input                                           std__pe3__lane5_strm0_data_valid  ;

  output                                          pe3__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane5_strm1_data_mask   ;
  input                                           std__pe3__lane5_strm1_data_valid  ;

  output                                          pe3__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane6_strm0_data_mask   ;
  input                                           std__pe3__lane6_strm0_data_valid  ;

  output                                          pe3__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane6_strm1_data_mask   ;
  input                                           std__pe3__lane6_strm1_data_valid  ;

  output                                          pe3__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane7_strm0_data_mask   ;
  input                                           std__pe3__lane7_strm0_data_valid  ;

  output                                          pe3__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane7_strm1_data_mask   ;
  input                                           std__pe3__lane7_strm1_data_valid  ;

  output                                          pe3__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane8_strm0_data_mask   ;
  input                                           std__pe3__lane8_strm0_data_valid  ;

  output                                          pe3__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane8_strm1_data_mask   ;
  input                                           std__pe3__lane8_strm1_data_valid  ;

  output                                          pe3__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane9_strm0_data_mask   ;
  input                                           std__pe3__lane9_strm0_data_valid  ;

  output                                          pe3__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane9_strm1_data_mask   ;
  input                                           std__pe3__lane9_strm1_data_valid  ;

  output                                          pe3__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane10_strm0_data_mask   ;
  input                                           std__pe3__lane10_strm0_data_valid  ;

  output                                          pe3__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane10_strm1_data_mask   ;
  input                                           std__pe3__lane10_strm1_data_valid  ;

  output                                          pe3__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane11_strm0_data_mask   ;
  input                                           std__pe3__lane11_strm0_data_valid  ;

  output                                          pe3__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane11_strm1_data_mask   ;
  input                                           std__pe3__lane11_strm1_data_valid  ;

  output                                          pe3__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane12_strm0_data_mask   ;
  input                                           std__pe3__lane12_strm0_data_valid  ;

  output                                          pe3__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane12_strm1_data_mask   ;
  input                                           std__pe3__lane12_strm1_data_valid  ;

  output                                          pe3__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane13_strm0_data_mask   ;
  input                                           std__pe3__lane13_strm0_data_valid  ;

  output                                          pe3__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane13_strm1_data_mask   ;
  input                                           std__pe3__lane13_strm1_data_valid  ;

  output                                          pe3__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane14_strm0_data_mask   ;
  input                                           std__pe3__lane14_strm0_data_valid  ;

  output                                          pe3__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane14_strm1_data_mask   ;
  input                                           std__pe3__lane14_strm1_data_valid  ;

  output                                          pe3__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane15_strm0_data_mask   ;
  input                                           std__pe3__lane15_strm0_data_valid  ;

  output                                          pe3__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane15_strm1_data_mask   ;
  input                                           std__pe3__lane15_strm1_data_valid  ;

  output                                          pe3__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane16_strm0_data_mask   ;
  input                                           std__pe3__lane16_strm0_data_valid  ;

  output                                          pe3__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane16_strm1_data_mask   ;
  input                                           std__pe3__lane16_strm1_data_valid  ;

  output                                          pe3__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane17_strm0_data_mask   ;
  input                                           std__pe3__lane17_strm0_data_valid  ;

  output                                          pe3__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane17_strm1_data_mask   ;
  input                                           std__pe3__lane17_strm1_data_valid  ;

  output                                          pe3__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane18_strm0_data_mask   ;
  input                                           std__pe3__lane18_strm0_data_valid  ;

  output                                          pe3__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane18_strm1_data_mask   ;
  input                                           std__pe3__lane18_strm1_data_valid  ;

  output                                          pe3__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane19_strm0_data_mask   ;
  input                                           std__pe3__lane19_strm0_data_valid  ;

  output                                          pe3__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane19_strm1_data_mask   ;
  input                                           std__pe3__lane19_strm1_data_valid  ;

  output                                          pe3__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane20_strm0_data_mask   ;
  input                                           std__pe3__lane20_strm0_data_valid  ;

  output                                          pe3__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane20_strm1_data_mask   ;
  input                                           std__pe3__lane20_strm1_data_valid  ;

  output                                          pe3__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane21_strm0_data_mask   ;
  input                                           std__pe3__lane21_strm0_data_valid  ;

  output                                          pe3__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane21_strm1_data_mask   ;
  input                                           std__pe3__lane21_strm1_data_valid  ;

  output                                          pe3__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane22_strm0_data_mask   ;
  input                                           std__pe3__lane22_strm0_data_valid  ;

  output                                          pe3__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane22_strm1_data_mask   ;
  input                                           std__pe3__lane22_strm1_data_valid  ;

  output                                          pe3__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane23_strm0_data_mask   ;
  input                                           std__pe3__lane23_strm0_data_valid  ;

  output                                          pe3__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane23_strm1_data_mask   ;
  input                                           std__pe3__lane23_strm1_data_valid  ;

  output                                          pe3__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane24_strm0_data_mask   ;
  input                                           std__pe3__lane24_strm0_data_valid  ;

  output                                          pe3__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane24_strm1_data_mask   ;
  input                                           std__pe3__lane24_strm1_data_valid  ;

  output                                          pe3__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane25_strm0_data_mask   ;
  input                                           std__pe3__lane25_strm0_data_valid  ;

  output                                          pe3__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane25_strm1_data_mask   ;
  input                                           std__pe3__lane25_strm1_data_valid  ;

  output                                          pe3__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane26_strm0_data_mask   ;
  input                                           std__pe3__lane26_strm0_data_valid  ;

  output                                          pe3__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane26_strm1_data_mask   ;
  input                                           std__pe3__lane26_strm1_data_valid  ;

  output                                          pe3__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane27_strm0_data_mask   ;
  input                                           std__pe3__lane27_strm0_data_valid  ;

  output                                          pe3__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane27_strm1_data_mask   ;
  input                                           std__pe3__lane27_strm1_data_valid  ;

  output                                          pe3__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane28_strm0_data_mask   ;
  input                                           std__pe3__lane28_strm0_data_valid  ;

  output                                          pe3__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane28_strm1_data_mask   ;
  input                                           std__pe3__lane28_strm1_data_valid  ;

  output                                          pe3__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane29_strm0_data_mask   ;
  input                                           std__pe3__lane29_strm0_data_valid  ;

  output                                          pe3__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane29_strm1_data_mask   ;
  input                                           std__pe3__lane29_strm1_data_valid  ;

  output                                          pe3__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane30_strm0_data_mask   ;
  input                                           std__pe3__lane30_strm0_data_valid  ;

  output                                          pe3__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane30_strm1_data_mask   ;
  input                                           std__pe3__lane30_strm1_data_valid  ;

  output                                          pe3__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane31_strm0_data_mask   ;
  input                                           std__pe3__lane31_strm0_data_valid  ;

  output                                          pe3__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe3__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe3__lane31_strm1_data_mask   ;
  input                                           std__pe3__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe4__peId                ;
  input                                         sys__pe4__allSynchronized     ;
  output                                        pe4__sys__thisSynchronized    ;
  output                                        pe4__sys__ready               ;
  output                                        pe4__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe4__oob_cntl            ;
  input                                         std__pe4__oob_valid           ;
  output                                        pe4__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe4__oob_type            ;
  output                                          pe4__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane0_strm0_data_mask   ;
  input                                           std__pe4__lane0_strm0_data_valid  ;

  output                                          pe4__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane0_strm1_data_mask   ;
  input                                           std__pe4__lane0_strm1_data_valid  ;

  output                                          pe4__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane1_strm0_data_mask   ;
  input                                           std__pe4__lane1_strm0_data_valid  ;

  output                                          pe4__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane1_strm1_data_mask   ;
  input                                           std__pe4__lane1_strm1_data_valid  ;

  output                                          pe4__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane2_strm0_data_mask   ;
  input                                           std__pe4__lane2_strm0_data_valid  ;

  output                                          pe4__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane2_strm1_data_mask   ;
  input                                           std__pe4__lane2_strm1_data_valid  ;

  output                                          pe4__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane3_strm0_data_mask   ;
  input                                           std__pe4__lane3_strm0_data_valid  ;

  output                                          pe4__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane3_strm1_data_mask   ;
  input                                           std__pe4__lane3_strm1_data_valid  ;

  output                                          pe4__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane4_strm0_data_mask   ;
  input                                           std__pe4__lane4_strm0_data_valid  ;

  output                                          pe4__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane4_strm1_data_mask   ;
  input                                           std__pe4__lane4_strm1_data_valid  ;

  output                                          pe4__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane5_strm0_data_mask   ;
  input                                           std__pe4__lane5_strm0_data_valid  ;

  output                                          pe4__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane5_strm1_data_mask   ;
  input                                           std__pe4__lane5_strm1_data_valid  ;

  output                                          pe4__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane6_strm0_data_mask   ;
  input                                           std__pe4__lane6_strm0_data_valid  ;

  output                                          pe4__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane6_strm1_data_mask   ;
  input                                           std__pe4__lane6_strm1_data_valid  ;

  output                                          pe4__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane7_strm0_data_mask   ;
  input                                           std__pe4__lane7_strm0_data_valid  ;

  output                                          pe4__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane7_strm1_data_mask   ;
  input                                           std__pe4__lane7_strm1_data_valid  ;

  output                                          pe4__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane8_strm0_data_mask   ;
  input                                           std__pe4__lane8_strm0_data_valid  ;

  output                                          pe4__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane8_strm1_data_mask   ;
  input                                           std__pe4__lane8_strm1_data_valid  ;

  output                                          pe4__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane9_strm0_data_mask   ;
  input                                           std__pe4__lane9_strm0_data_valid  ;

  output                                          pe4__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane9_strm1_data_mask   ;
  input                                           std__pe4__lane9_strm1_data_valid  ;

  output                                          pe4__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane10_strm0_data_mask   ;
  input                                           std__pe4__lane10_strm0_data_valid  ;

  output                                          pe4__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane10_strm1_data_mask   ;
  input                                           std__pe4__lane10_strm1_data_valid  ;

  output                                          pe4__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane11_strm0_data_mask   ;
  input                                           std__pe4__lane11_strm0_data_valid  ;

  output                                          pe4__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane11_strm1_data_mask   ;
  input                                           std__pe4__lane11_strm1_data_valid  ;

  output                                          pe4__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane12_strm0_data_mask   ;
  input                                           std__pe4__lane12_strm0_data_valid  ;

  output                                          pe4__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane12_strm1_data_mask   ;
  input                                           std__pe4__lane12_strm1_data_valid  ;

  output                                          pe4__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane13_strm0_data_mask   ;
  input                                           std__pe4__lane13_strm0_data_valid  ;

  output                                          pe4__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane13_strm1_data_mask   ;
  input                                           std__pe4__lane13_strm1_data_valid  ;

  output                                          pe4__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane14_strm0_data_mask   ;
  input                                           std__pe4__lane14_strm0_data_valid  ;

  output                                          pe4__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane14_strm1_data_mask   ;
  input                                           std__pe4__lane14_strm1_data_valid  ;

  output                                          pe4__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane15_strm0_data_mask   ;
  input                                           std__pe4__lane15_strm0_data_valid  ;

  output                                          pe4__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane15_strm1_data_mask   ;
  input                                           std__pe4__lane15_strm1_data_valid  ;

  output                                          pe4__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane16_strm0_data_mask   ;
  input                                           std__pe4__lane16_strm0_data_valid  ;

  output                                          pe4__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane16_strm1_data_mask   ;
  input                                           std__pe4__lane16_strm1_data_valid  ;

  output                                          pe4__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane17_strm0_data_mask   ;
  input                                           std__pe4__lane17_strm0_data_valid  ;

  output                                          pe4__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane17_strm1_data_mask   ;
  input                                           std__pe4__lane17_strm1_data_valid  ;

  output                                          pe4__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane18_strm0_data_mask   ;
  input                                           std__pe4__lane18_strm0_data_valid  ;

  output                                          pe4__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane18_strm1_data_mask   ;
  input                                           std__pe4__lane18_strm1_data_valid  ;

  output                                          pe4__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane19_strm0_data_mask   ;
  input                                           std__pe4__lane19_strm0_data_valid  ;

  output                                          pe4__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane19_strm1_data_mask   ;
  input                                           std__pe4__lane19_strm1_data_valid  ;

  output                                          pe4__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane20_strm0_data_mask   ;
  input                                           std__pe4__lane20_strm0_data_valid  ;

  output                                          pe4__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane20_strm1_data_mask   ;
  input                                           std__pe4__lane20_strm1_data_valid  ;

  output                                          pe4__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane21_strm0_data_mask   ;
  input                                           std__pe4__lane21_strm0_data_valid  ;

  output                                          pe4__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane21_strm1_data_mask   ;
  input                                           std__pe4__lane21_strm1_data_valid  ;

  output                                          pe4__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane22_strm0_data_mask   ;
  input                                           std__pe4__lane22_strm0_data_valid  ;

  output                                          pe4__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane22_strm1_data_mask   ;
  input                                           std__pe4__lane22_strm1_data_valid  ;

  output                                          pe4__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane23_strm0_data_mask   ;
  input                                           std__pe4__lane23_strm0_data_valid  ;

  output                                          pe4__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane23_strm1_data_mask   ;
  input                                           std__pe4__lane23_strm1_data_valid  ;

  output                                          pe4__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane24_strm0_data_mask   ;
  input                                           std__pe4__lane24_strm0_data_valid  ;

  output                                          pe4__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane24_strm1_data_mask   ;
  input                                           std__pe4__lane24_strm1_data_valid  ;

  output                                          pe4__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane25_strm0_data_mask   ;
  input                                           std__pe4__lane25_strm0_data_valid  ;

  output                                          pe4__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane25_strm1_data_mask   ;
  input                                           std__pe4__lane25_strm1_data_valid  ;

  output                                          pe4__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane26_strm0_data_mask   ;
  input                                           std__pe4__lane26_strm0_data_valid  ;

  output                                          pe4__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane26_strm1_data_mask   ;
  input                                           std__pe4__lane26_strm1_data_valid  ;

  output                                          pe4__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane27_strm0_data_mask   ;
  input                                           std__pe4__lane27_strm0_data_valid  ;

  output                                          pe4__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane27_strm1_data_mask   ;
  input                                           std__pe4__lane27_strm1_data_valid  ;

  output                                          pe4__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane28_strm0_data_mask   ;
  input                                           std__pe4__lane28_strm0_data_valid  ;

  output                                          pe4__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane28_strm1_data_mask   ;
  input                                           std__pe4__lane28_strm1_data_valid  ;

  output                                          pe4__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane29_strm0_data_mask   ;
  input                                           std__pe4__lane29_strm0_data_valid  ;

  output                                          pe4__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane29_strm1_data_mask   ;
  input                                           std__pe4__lane29_strm1_data_valid  ;

  output                                          pe4__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane30_strm0_data_mask   ;
  input                                           std__pe4__lane30_strm0_data_valid  ;

  output                                          pe4__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane30_strm1_data_mask   ;
  input                                           std__pe4__lane30_strm1_data_valid  ;

  output                                          pe4__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane31_strm0_data_mask   ;
  input                                           std__pe4__lane31_strm0_data_valid  ;

  output                                          pe4__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe4__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe4__lane31_strm1_data_mask   ;
  input                                           std__pe4__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe5__peId                ;
  input                                         sys__pe5__allSynchronized     ;
  output                                        pe5__sys__thisSynchronized    ;
  output                                        pe5__sys__ready               ;
  output                                        pe5__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe5__oob_cntl            ;
  input                                         std__pe5__oob_valid           ;
  output                                        pe5__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe5__oob_type            ;
  output                                          pe5__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane0_strm0_data_mask   ;
  input                                           std__pe5__lane0_strm0_data_valid  ;

  output                                          pe5__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane0_strm1_data_mask   ;
  input                                           std__pe5__lane0_strm1_data_valid  ;

  output                                          pe5__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane1_strm0_data_mask   ;
  input                                           std__pe5__lane1_strm0_data_valid  ;

  output                                          pe5__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane1_strm1_data_mask   ;
  input                                           std__pe5__lane1_strm1_data_valid  ;

  output                                          pe5__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane2_strm0_data_mask   ;
  input                                           std__pe5__lane2_strm0_data_valid  ;

  output                                          pe5__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane2_strm1_data_mask   ;
  input                                           std__pe5__lane2_strm1_data_valid  ;

  output                                          pe5__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane3_strm0_data_mask   ;
  input                                           std__pe5__lane3_strm0_data_valid  ;

  output                                          pe5__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane3_strm1_data_mask   ;
  input                                           std__pe5__lane3_strm1_data_valid  ;

  output                                          pe5__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane4_strm0_data_mask   ;
  input                                           std__pe5__lane4_strm0_data_valid  ;

  output                                          pe5__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane4_strm1_data_mask   ;
  input                                           std__pe5__lane4_strm1_data_valid  ;

  output                                          pe5__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane5_strm0_data_mask   ;
  input                                           std__pe5__lane5_strm0_data_valid  ;

  output                                          pe5__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane5_strm1_data_mask   ;
  input                                           std__pe5__lane5_strm1_data_valid  ;

  output                                          pe5__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane6_strm0_data_mask   ;
  input                                           std__pe5__lane6_strm0_data_valid  ;

  output                                          pe5__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane6_strm1_data_mask   ;
  input                                           std__pe5__lane6_strm1_data_valid  ;

  output                                          pe5__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane7_strm0_data_mask   ;
  input                                           std__pe5__lane7_strm0_data_valid  ;

  output                                          pe5__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane7_strm1_data_mask   ;
  input                                           std__pe5__lane7_strm1_data_valid  ;

  output                                          pe5__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane8_strm0_data_mask   ;
  input                                           std__pe5__lane8_strm0_data_valid  ;

  output                                          pe5__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane8_strm1_data_mask   ;
  input                                           std__pe5__lane8_strm1_data_valid  ;

  output                                          pe5__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane9_strm0_data_mask   ;
  input                                           std__pe5__lane9_strm0_data_valid  ;

  output                                          pe5__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane9_strm1_data_mask   ;
  input                                           std__pe5__lane9_strm1_data_valid  ;

  output                                          pe5__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane10_strm0_data_mask   ;
  input                                           std__pe5__lane10_strm0_data_valid  ;

  output                                          pe5__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane10_strm1_data_mask   ;
  input                                           std__pe5__lane10_strm1_data_valid  ;

  output                                          pe5__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane11_strm0_data_mask   ;
  input                                           std__pe5__lane11_strm0_data_valid  ;

  output                                          pe5__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane11_strm1_data_mask   ;
  input                                           std__pe5__lane11_strm1_data_valid  ;

  output                                          pe5__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane12_strm0_data_mask   ;
  input                                           std__pe5__lane12_strm0_data_valid  ;

  output                                          pe5__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane12_strm1_data_mask   ;
  input                                           std__pe5__lane12_strm1_data_valid  ;

  output                                          pe5__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane13_strm0_data_mask   ;
  input                                           std__pe5__lane13_strm0_data_valid  ;

  output                                          pe5__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane13_strm1_data_mask   ;
  input                                           std__pe5__lane13_strm1_data_valid  ;

  output                                          pe5__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane14_strm0_data_mask   ;
  input                                           std__pe5__lane14_strm0_data_valid  ;

  output                                          pe5__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane14_strm1_data_mask   ;
  input                                           std__pe5__lane14_strm1_data_valid  ;

  output                                          pe5__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane15_strm0_data_mask   ;
  input                                           std__pe5__lane15_strm0_data_valid  ;

  output                                          pe5__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane15_strm1_data_mask   ;
  input                                           std__pe5__lane15_strm1_data_valid  ;

  output                                          pe5__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane16_strm0_data_mask   ;
  input                                           std__pe5__lane16_strm0_data_valid  ;

  output                                          pe5__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane16_strm1_data_mask   ;
  input                                           std__pe5__lane16_strm1_data_valid  ;

  output                                          pe5__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane17_strm0_data_mask   ;
  input                                           std__pe5__lane17_strm0_data_valid  ;

  output                                          pe5__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane17_strm1_data_mask   ;
  input                                           std__pe5__lane17_strm1_data_valid  ;

  output                                          pe5__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane18_strm0_data_mask   ;
  input                                           std__pe5__lane18_strm0_data_valid  ;

  output                                          pe5__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane18_strm1_data_mask   ;
  input                                           std__pe5__lane18_strm1_data_valid  ;

  output                                          pe5__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane19_strm0_data_mask   ;
  input                                           std__pe5__lane19_strm0_data_valid  ;

  output                                          pe5__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane19_strm1_data_mask   ;
  input                                           std__pe5__lane19_strm1_data_valid  ;

  output                                          pe5__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane20_strm0_data_mask   ;
  input                                           std__pe5__lane20_strm0_data_valid  ;

  output                                          pe5__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane20_strm1_data_mask   ;
  input                                           std__pe5__lane20_strm1_data_valid  ;

  output                                          pe5__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane21_strm0_data_mask   ;
  input                                           std__pe5__lane21_strm0_data_valid  ;

  output                                          pe5__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane21_strm1_data_mask   ;
  input                                           std__pe5__lane21_strm1_data_valid  ;

  output                                          pe5__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane22_strm0_data_mask   ;
  input                                           std__pe5__lane22_strm0_data_valid  ;

  output                                          pe5__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane22_strm1_data_mask   ;
  input                                           std__pe5__lane22_strm1_data_valid  ;

  output                                          pe5__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane23_strm0_data_mask   ;
  input                                           std__pe5__lane23_strm0_data_valid  ;

  output                                          pe5__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane23_strm1_data_mask   ;
  input                                           std__pe5__lane23_strm1_data_valid  ;

  output                                          pe5__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane24_strm0_data_mask   ;
  input                                           std__pe5__lane24_strm0_data_valid  ;

  output                                          pe5__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane24_strm1_data_mask   ;
  input                                           std__pe5__lane24_strm1_data_valid  ;

  output                                          pe5__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane25_strm0_data_mask   ;
  input                                           std__pe5__lane25_strm0_data_valid  ;

  output                                          pe5__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane25_strm1_data_mask   ;
  input                                           std__pe5__lane25_strm1_data_valid  ;

  output                                          pe5__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane26_strm0_data_mask   ;
  input                                           std__pe5__lane26_strm0_data_valid  ;

  output                                          pe5__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane26_strm1_data_mask   ;
  input                                           std__pe5__lane26_strm1_data_valid  ;

  output                                          pe5__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane27_strm0_data_mask   ;
  input                                           std__pe5__lane27_strm0_data_valid  ;

  output                                          pe5__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane27_strm1_data_mask   ;
  input                                           std__pe5__lane27_strm1_data_valid  ;

  output                                          pe5__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane28_strm0_data_mask   ;
  input                                           std__pe5__lane28_strm0_data_valid  ;

  output                                          pe5__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane28_strm1_data_mask   ;
  input                                           std__pe5__lane28_strm1_data_valid  ;

  output                                          pe5__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane29_strm0_data_mask   ;
  input                                           std__pe5__lane29_strm0_data_valid  ;

  output                                          pe5__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane29_strm1_data_mask   ;
  input                                           std__pe5__lane29_strm1_data_valid  ;

  output                                          pe5__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane30_strm0_data_mask   ;
  input                                           std__pe5__lane30_strm0_data_valid  ;

  output                                          pe5__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane30_strm1_data_mask   ;
  input                                           std__pe5__lane30_strm1_data_valid  ;

  output                                          pe5__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane31_strm0_data_mask   ;
  input                                           std__pe5__lane31_strm0_data_valid  ;

  output                                          pe5__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe5__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe5__lane31_strm1_data_mask   ;
  input                                           std__pe5__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe6__peId                ;
  input                                         sys__pe6__allSynchronized     ;
  output                                        pe6__sys__thisSynchronized    ;
  output                                        pe6__sys__ready               ;
  output                                        pe6__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe6__oob_cntl            ;
  input                                         std__pe6__oob_valid           ;
  output                                        pe6__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe6__oob_type            ;
  output                                          pe6__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane0_strm0_data_mask   ;
  input                                           std__pe6__lane0_strm0_data_valid  ;

  output                                          pe6__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane0_strm1_data_mask   ;
  input                                           std__pe6__lane0_strm1_data_valid  ;

  output                                          pe6__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane1_strm0_data_mask   ;
  input                                           std__pe6__lane1_strm0_data_valid  ;

  output                                          pe6__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane1_strm1_data_mask   ;
  input                                           std__pe6__lane1_strm1_data_valid  ;

  output                                          pe6__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane2_strm0_data_mask   ;
  input                                           std__pe6__lane2_strm0_data_valid  ;

  output                                          pe6__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane2_strm1_data_mask   ;
  input                                           std__pe6__lane2_strm1_data_valid  ;

  output                                          pe6__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane3_strm0_data_mask   ;
  input                                           std__pe6__lane3_strm0_data_valid  ;

  output                                          pe6__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane3_strm1_data_mask   ;
  input                                           std__pe6__lane3_strm1_data_valid  ;

  output                                          pe6__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane4_strm0_data_mask   ;
  input                                           std__pe6__lane4_strm0_data_valid  ;

  output                                          pe6__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane4_strm1_data_mask   ;
  input                                           std__pe6__lane4_strm1_data_valid  ;

  output                                          pe6__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane5_strm0_data_mask   ;
  input                                           std__pe6__lane5_strm0_data_valid  ;

  output                                          pe6__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane5_strm1_data_mask   ;
  input                                           std__pe6__lane5_strm1_data_valid  ;

  output                                          pe6__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane6_strm0_data_mask   ;
  input                                           std__pe6__lane6_strm0_data_valid  ;

  output                                          pe6__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane6_strm1_data_mask   ;
  input                                           std__pe6__lane6_strm1_data_valid  ;

  output                                          pe6__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane7_strm0_data_mask   ;
  input                                           std__pe6__lane7_strm0_data_valid  ;

  output                                          pe6__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane7_strm1_data_mask   ;
  input                                           std__pe6__lane7_strm1_data_valid  ;

  output                                          pe6__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane8_strm0_data_mask   ;
  input                                           std__pe6__lane8_strm0_data_valid  ;

  output                                          pe6__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane8_strm1_data_mask   ;
  input                                           std__pe6__lane8_strm1_data_valid  ;

  output                                          pe6__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane9_strm0_data_mask   ;
  input                                           std__pe6__lane9_strm0_data_valid  ;

  output                                          pe6__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane9_strm1_data_mask   ;
  input                                           std__pe6__lane9_strm1_data_valid  ;

  output                                          pe6__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane10_strm0_data_mask   ;
  input                                           std__pe6__lane10_strm0_data_valid  ;

  output                                          pe6__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane10_strm1_data_mask   ;
  input                                           std__pe6__lane10_strm1_data_valid  ;

  output                                          pe6__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane11_strm0_data_mask   ;
  input                                           std__pe6__lane11_strm0_data_valid  ;

  output                                          pe6__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane11_strm1_data_mask   ;
  input                                           std__pe6__lane11_strm1_data_valid  ;

  output                                          pe6__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane12_strm0_data_mask   ;
  input                                           std__pe6__lane12_strm0_data_valid  ;

  output                                          pe6__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane12_strm1_data_mask   ;
  input                                           std__pe6__lane12_strm1_data_valid  ;

  output                                          pe6__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane13_strm0_data_mask   ;
  input                                           std__pe6__lane13_strm0_data_valid  ;

  output                                          pe6__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane13_strm1_data_mask   ;
  input                                           std__pe6__lane13_strm1_data_valid  ;

  output                                          pe6__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane14_strm0_data_mask   ;
  input                                           std__pe6__lane14_strm0_data_valid  ;

  output                                          pe6__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane14_strm1_data_mask   ;
  input                                           std__pe6__lane14_strm1_data_valid  ;

  output                                          pe6__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane15_strm0_data_mask   ;
  input                                           std__pe6__lane15_strm0_data_valid  ;

  output                                          pe6__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane15_strm1_data_mask   ;
  input                                           std__pe6__lane15_strm1_data_valid  ;

  output                                          pe6__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane16_strm0_data_mask   ;
  input                                           std__pe6__lane16_strm0_data_valid  ;

  output                                          pe6__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane16_strm1_data_mask   ;
  input                                           std__pe6__lane16_strm1_data_valid  ;

  output                                          pe6__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane17_strm0_data_mask   ;
  input                                           std__pe6__lane17_strm0_data_valid  ;

  output                                          pe6__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane17_strm1_data_mask   ;
  input                                           std__pe6__lane17_strm1_data_valid  ;

  output                                          pe6__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane18_strm0_data_mask   ;
  input                                           std__pe6__lane18_strm0_data_valid  ;

  output                                          pe6__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane18_strm1_data_mask   ;
  input                                           std__pe6__lane18_strm1_data_valid  ;

  output                                          pe6__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane19_strm0_data_mask   ;
  input                                           std__pe6__lane19_strm0_data_valid  ;

  output                                          pe6__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane19_strm1_data_mask   ;
  input                                           std__pe6__lane19_strm1_data_valid  ;

  output                                          pe6__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane20_strm0_data_mask   ;
  input                                           std__pe6__lane20_strm0_data_valid  ;

  output                                          pe6__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane20_strm1_data_mask   ;
  input                                           std__pe6__lane20_strm1_data_valid  ;

  output                                          pe6__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane21_strm0_data_mask   ;
  input                                           std__pe6__lane21_strm0_data_valid  ;

  output                                          pe6__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane21_strm1_data_mask   ;
  input                                           std__pe6__lane21_strm1_data_valid  ;

  output                                          pe6__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane22_strm0_data_mask   ;
  input                                           std__pe6__lane22_strm0_data_valid  ;

  output                                          pe6__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane22_strm1_data_mask   ;
  input                                           std__pe6__lane22_strm1_data_valid  ;

  output                                          pe6__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane23_strm0_data_mask   ;
  input                                           std__pe6__lane23_strm0_data_valid  ;

  output                                          pe6__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane23_strm1_data_mask   ;
  input                                           std__pe6__lane23_strm1_data_valid  ;

  output                                          pe6__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane24_strm0_data_mask   ;
  input                                           std__pe6__lane24_strm0_data_valid  ;

  output                                          pe6__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane24_strm1_data_mask   ;
  input                                           std__pe6__lane24_strm1_data_valid  ;

  output                                          pe6__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane25_strm0_data_mask   ;
  input                                           std__pe6__lane25_strm0_data_valid  ;

  output                                          pe6__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane25_strm1_data_mask   ;
  input                                           std__pe6__lane25_strm1_data_valid  ;

  output                                          pe6__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane26_strm0_data_mask   ;
  input                                           std__pe6__lane26_strm0_data_valid  ;

  output                                          pe6__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane26_strm1_data_mask   ;
  input                                           std__pe6__lane26_strm1_data_valid  ;

  output                                          pe6__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane27_strm0_data_mask   ;
  input                                           std__pe6__lane27_strm0_data_valid  ;

  output                                          pe6__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane27_strm1_data_mask   ;
  input                                           std__pe6__lane27_strm1_data_valid  ;

  output                                          pe6__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane28_strm0_data_mask   ;
  input                                           std__pe6__lane28_strm0_data_valid  ;

  output                                          pe6__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane28_strm1_data_mask   ;
  input                                           std__pe6__lane28_strm1_data_valid  ;

  output                                          pe6__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane29_strm0_data_mask   ;
  input                                           std__pe6__lane29_strm0_data_valid  ;

  output                                          pe6__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane29_strm1_data_mask   ;
  input                                           std__pe6__lane29_strm1_data_valid  ;

  output                                          pe6__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane30_strm0_data_mask   ;
  input                                           std__pe6__lane30_strm0_data_valid  ;

  output                                          pe6__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane30_strm1_data_mask   ;
  input                                           std__pe6__lane30_strm1_data_valid  ;

  output                                          pe6__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane31_strm0_data_mask   ;
  input                                           std__pe6__lane31_strm0_data_valid  ;

  output                                          pe6__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe6__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe6__lane31_strm1_data_mask   ;
  input                                           std__pe6__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe7__peId                ;
  input                                         sys__pe7__allSynchronized     ;
  output                                        pe7__sys__thisSynchronized    ;
  output                                        pe7__sys__ready               ;
  output                                        pe7__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe7__oob_cntl            ;
  input                                         std__pe7__oob_valid           ;
  output                                        pe7__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe7__oob_type            ;
  output                                          pe7__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane0_strm0_data_mask   ;
  input                                           std__pe7__lane0_strm0_data_valid  ;

  output                                          pe7__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane0_strm1_data_mask   ;
  input                                           std__pe7__lane0_strm1_data_valid  ;

  output                                          pe7__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane1_strm0_data_mask   ;
  input                                           std__pe7__lane1_strm0_data_valid  ;

  output                                          pe7__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane1_strm1_data_mask   ;
  input                                           std__pe7__lane1_strm1_data_valid  ;

  output                                          pe7__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane2_strm0_data_mask   ;
  input                                           std__pe7__lane2_strm0_data_valid  ;

  output                                          pe7__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane2_strm1_data_mask   ;
  input                                           std__pe7__lane2_strm1_data_valid  ;

  output                                          pe7__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane3_strm0_data_mask   ;
  input                                           std__pe7__lane3_strm0_data_valid  ;

  output                                          pe7__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane3_strm1_data_mask   ;
  input                                           std__pe7__lane3_strm1_data_valid  ;

  output                                          pe7__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane4_strm0_data_mask   ;
  input                                           std__pe7__lane4_strm0_data_valid  ;

  output                                          pe7__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane4_strm1_data_mask   ;
  input                                           std__pe7__lane4_strm1_data_valid  ;

  output                                          pe7__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane5_strm0_data_mask   ;
  input                                           std__pe7__lane5_strm0_data_valid  ;

  output                                          pe7__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane5_strm1_data_mask   ;
  input                                           std__pe7__lane5_strm1_data_valid  ;

  output                                          pe7__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane6_strm0_data_mask   ;
  input                                           std__pe7__lane6_strm0_data_valid  ;

  output                                          pe7__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane6_strm1_data_mask   ;
  input                                           std__pe7__lane6_strm1_data_valid  ;

  output                                          pe7__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane7_strm0_data_mask   ;
  input                                           std__pe7__lane7_strm0_data_valid  ;

  output                                          pe7__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane7_strm1_data_mask   ;
  input                                           std__pe7__lane7_strm1_data_valid  ;

  output                                          pe7__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane8_strm0_data_mask   ;
  input                                           std__pe7__lane8_strm0_data_valid  ;

  output                                          pe7__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane8_strm1_data_mask   ;
  input                                           std__pe7__lane8_strm1_data_valid  ;

  output                                          pe7__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane9_strm0_data_mask   ;
  input                                           std__pe7__lane9_strm0_data_valid  ;

  output                                          pe7__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane9_strm1_data_mask   ;
  input                                           std__pe7__lane9_strm1_data_valid  ;

  output                                          pe7__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane10_strm0_data_mask   ;
  input                                           std__pe7__lane10_strm0_data_valid  ;

  output                                          pe7__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane10_strm1_data_mask   ;
  input                                           std__pe7__lane10_strm1_data_valid  ;

  output                                          pe7__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane11_strm0_data_mask   ;
  input                                           std__pe7__lane11_strm0_data_valid  ;

  output                                          pe7__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane11_strm1_data_mask   ;
  input                                           std__pe7__lane11_strm1_data_valid  ;

  output                                          pe7__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane12_strm0_data_mask   ;
  input                                           std__pe7__lane12_strm0_data_valid  ;

  output                                          pe7__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane12_strm1_data_mask   ;
  input                                           std__pe7__lane12_strm1_data_valid  ;

  output                                          pe7__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane13_strm0_data_mask   ;
  input                                           std__pe7__lane13_strm0_data_valid  ;

  output                                          pe7__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane13_strm1_data_mask   ;
  input                                           std__pe7__lane13_strm1_data_valid  ;

  output                                          pe7__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane14_strm0_data_mask   ;
  input                                           std__pe7__lane14_strm0_data_valid  ;

  output                                          pe7__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane14_strm1_data_mask   ;
  input                                           std__pe7__lane14_strm1_data_valid  ;

  output                                          pe7__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane15_strm0_data_mask   ;
  input                                           std__pe7__lane15_strm0_data_valid  ;

  output                                          pe7__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane15_strm1_data_mask   ;
  input                                           std__pe7__lane15_strm1_data_valid  ;

  output                                          pe7__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane16_strm0_data_mask   ;
  input                                           std__pe7__lane16_strm0_data_valid  ;

  output                                          pe7__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane16_strm1_data_mask   ;
  input                                           std__pe7__lane16_strm1_data_valid  ;

  output                                          pe7__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane17_strm0_data_mask   ;
  input                                           std__pe7__lane17_strm0_data_valid  ;

  output                                          pe7__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane17_strm1_data_mask   ;
  input                                           std__pe7__lane17_strm1_data_valid  ;

  output                                          pe7__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane18_strm0_data_mask   ;
  input                                           std__pe7__lane18_strm0_data_valid  ;

  output                                          pe7__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane18_strm1_data_mask   ;
  input                                           std__pe7__lane18_strm1_data_valid  ;

  output                                          pe7__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane19_strm0_data_mask   ;
  input                                           std__pe7__lane19_strm0_data_valid  ;

  output                                          pe7__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane19_strm1_data_mask   ;
  input                                           std__pe7__lane19_strm1_data_valid  ;

  output                                          pe7__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane20_strm0_data_mask   ;
  input                                           std__pe7__lane20_strm0_data_valid  ;

  output                                          pe7__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane20_strm1_data_mask   ;
  input                                           std__pe7__lane20_strm1_data_valid  ;

  output                                          pe7__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane21_strm0_data_mask   ;
  input                                           std__pe7__lane21_strm0_data_valid  ;

  output                                          pe7__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane21_strm1_data_mask   ;
  input                                           std__pe7__lane21_strm1_data_valid  ;

  output                                          pe7__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane22_strm0_data_mask   ;
  input                                           std__pe7__lane22_strm0_data_valid  ;

  output                                          pe7__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane22_strm1_data_mask   ;
  input                                           std__pe7__lane22_strm1_data_valid  ;

  output                                          pe7__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane23_strm0_data_mask   ;
  input                                           std__pe7__lane23_strm0_data_valid  ;

  output                                          pe7__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane23_strm1_data_mask   ;
  input                                           std__pe7__lane23_strm1_data_valid  ;

  output                                          pe7__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane24_strm0_data_mask   ;
  input                                           std__pe7__lane24_strm0_data_valid  ;

  output                                          pe7__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane24_strm1_data_mask   ;
  input                                           std__pe7__lane24_strm1_data_valid  ;

  output                                          pe7__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane25_strm0_data_mask   ;
  input                                           std__pe7__lane25_strm0_data_valid  ;

  output                                          pe7__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane25_strm1_data_mask   ;
  input                                           std__pe7__lane25_strm1_data_valid  ;

  output                                          pe7__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane26_strm0_data_mask   ;
  input                                           std__pe7__lane26_strm0_data_valid  ;

  output                                          pe7__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane26_strm1_data_mask   ;
  input                                           std__pe7__lane26_strm1_data_valid  ;

  output                                          pe7__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane27_strm0_data_mask   ;
  input                                           std__pe7__lane27_strm0_data_valid  ;

  output                                          pe7__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane27_strm1_data_mask   ;
  input                                           std__pe7__lane27_strm1_data_valid  ;

  output                                          pe7__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane28_strm0_data_mask   ;
  input                                           std__pe7__lane28_strm0_data_valid  ;

  output                                          pe7__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane28_strm1_data_mask   ;
  input                                           std__pe7__lane28_strm1_data_valid  ;

  output                                          pe7__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane29_strm0_data_mask   ;
  input                                           std__pe7__lane29_strm0_data_valid  ;

  output                                          pe7__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane29_strm1_data_mask   ;
  input                                           std__pe7__lane29_strm1_data_valid  ;

  output                                          pe7__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane30_strm0_data_mask   ;
  input                                           std__pe7__lane30_strm0_data_valid  ;

  output                                          pe7__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane30_strm1_data_mask   ;
  input                                           std__pe7__lane30_strm1_data_valid  ;

  output                                          pe7__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane31_strm0_data_mask   ;
  input                                           std__pe7__lane31_strm0_data_valid  ;

  output                                          pe7__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe7__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe7__lane31_strm1_data_mask   ;
  input                                           std__pe7__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe8__peId                ;
  input                                         sys__pe8__allSynchronized     ;
  output                                        pe8__sys__thisSynchronized    ;
  output                                        pe8__sys__ready               ;
  output                                        pe8__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe8__oob_cntl            ;
  input                                         std__pe8__oob_valid           ;
  output                                        pe8__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe8__oob_type            ;
  output                                          pe8__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane0_strm0_data_mask   ;
  input                                           std__pe8__lane0_strm0_data_valid  ;

  output                                          pe8__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane0_strm1_data_mask   ;
  input                                           std__pe8__lane0_strm1_data_valid  ;

  output                                          pe8__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane1_strm0_data_mask   ;
  input                                           std__pe8__lane1_strm0_data_valid  ;

  output                                          pe8__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane1_strm1_data_mask   ;
  input                                           std__pe8__lane1_strm1_data_valid  ;

  output                                          pe8__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane2_strm0_data_mask   ;
  input                                           std__pe8__lane2_strm0_data_valid  ;

  output                                          pe8__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane2_strm1_data_mask   ;
  input                                           std__pe8__lane2_strm1_data_valid  ;

  output                                          pe8__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane3_strm0_data_mask   ;
  input                                           std__pe8__lane3_strm0_data_valid  ;

  output                                          pe8__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane3_strm1_data_mask   ;
  input                                           std__pe8__lane3_strm1_data_valid  ;

  output                                          pe8__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane4_strm0_data_mask   ;
  input                                           std__pe8__lane4_strm0_data_valid  ;

  output                                          pe8__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane4_strm1_data_mask   ;
  input                                           std__pe8__lane4_strm1_data_valid  ;

  output                                          pe8__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane5_strm0_data_mask   ;
  input                                           std__pe8__lane5_strm0_data_valid  ;

  output                                          pe8__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane5_strm1_data_mask   ;
  input                                           std__pe8__lane5_strm1_data_valid  ;

  output                                          pe8__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane6_strm0_data_mask   ;
  input                                           std__pe8__lane6_strm0_data_valid  ;

  output                                          pe8__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane6_strm1_data_mask   ;
  input                                           std__pe8__lane6_strm1_data_valid  ;

  output                                          pe8__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane7_strm0_data_mask   ;
  input                                           std__pe8__lane7_strm0_data_valid  ;

  output                                          pe8__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane7_strm1_data_mask   ;
  input                                           std__pe8__lane7_strm1_data_valid  ;

  output                                          pe8__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane8_strm0_data_mask   ;
  input                                           std__pe8__lane8_strm0_data_valid  ;

  output                                          pe8__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane8_strm1_data_mask   ;
  input                                           std__pe8__lane8_strm1_data_valid  ;

  output                                          pe8__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane9_strm0_data_mask   ;
  input                                           std__pe8__lane9_strm0_data_valid  ;

  output                                          pe8__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane9_strm1_data_mask   ;
  input                                           std__pe8__lane9_strm1_data_valid  ;

  output                                          pe8__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane10_strm0_data_mask   ;
  input                                           std__pe8__lane10_strm0_data_valid  ;

  output                                          pe8__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane10_strm1_data_mask   ;
  input                                           std__pe8__lane10_strm1_data_valid  ;

  output                                          pe8__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane11_strm0_data_mask   ;
  input                                           std__pe8__lane11_strm0_data_valid  ;

  output                                          pe8__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane11_strm1_data_mask   ;
  input                                           std__pe8__lane11_strm1_data_valid  ;

  output                                          pe8__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane12_strm0_data_mask   ;
  input                                           std__pe8__lane12_strm0_data_valid  ;

  output                                          pe8__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane12_strm1_data_mask   ;
  input                                           std__pe8__lane12_strm1_data_valid  ;

  output                                          pe8__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane13_strm0_data_mask   ;
  input                                           std__pe8__lane13_strm0_data_valid  ;

  output                                          pe8__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane13_strm1_data_mask   ;
  input                                           std__pe8__lane13_strm1_data_valid  ;

  output                                          pe8__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane14_strm0_data_mask   ;
  input                                           std__pe8__lane14_strm0_data_valid  ;

  output                                          pe8__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane14_strm1_data_mask   ;
  input                                           std__pe8__lane14_strm1_data_valid  ;

  output                                          pe8__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane15_strm0_data_mask   ;
  input                                           std__pe8__lane15_strm0_data_valid  ;

  output                                          pe8__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane15_strm1_data_mask   ;
  input                                           std__pe8__lane15_strm1_data_valid  ;

  output                                          pe8__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane16_strm0_data_mask   ;
  input                                           std__pe8__lane16_strm0_data_valid  ;

  output                                          pe8__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane16_strm1_data_mask   ;
  input                                           std__pe8__lane16_strm1_data_valid  ;

  output                                          pe8__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane17_strm0_data_mask   ;
  input                                           std__pe8__lane17_strm0_data_valid  ;

  output                                          pe8__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane17_strm1_data_mask   ;
  input                                           std__pe8__lane17_strm1_data_valid  ;

  output                                          pe8__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane18_strm0_data_mask   ;
  input                                           std__pe8__lane18_strm0_data_valid  ;

  output                                          pe8__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane18_strm1_data_mask   ;
  input                                           std__pe8__lane18_strm1_data_valid  ;

  output                                          pe8__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane19_strm0_data_mask   ;
  input                                           std__pe8__lane19_strm0_data_valid  ;

  output                                          pe8__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane19_strm1_data_mask   ;
  input                                           std__pe8__lane19_strm1_data_valid  ;

  output                                          pe8__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane20_strm0_data_mask   ;
  input                                           std__pe8__lane20_strm0_data_valid  ;

  output                                          pe8__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane20_strm1_data_mask   ;
  input                                           std__pe8__lane20_strm1_data_valid  ;

  output                                          pe8__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane21_strm0_data_mask   ;
  input                                           std__pe8__lane21_strm0_data_valid  ;

  output                                          pe8__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane21_strm1_data_mask   ;
  input                                           std__pe8__lane21_strm1_data_valid  ;

  output                                          pe8__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane22_strm0_data_mask   ;
  input                                           std__pe8__lane22_strm0_data_valid  ;

  output                                          pe8__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane22_strm1_data_mask   ;
  input                                           std__pe8__lane22_strm1_data_valid  ;

  output                                          pe8__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane23_strm0_data_mask   ;
  input                                           std__pe8__lane23_strm0_data_valid  ;

  output                                          pe8__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane23_strm1_data_mask   ;
  input                                           std__pe8__lane23_strm1_data_valid  ;

  output                                          pe8__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane24_strm0_data_mask   ;
  input                                           std__pe8__lane24_strm0_data_valid  ;

  output                                          pe8__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane24_strm1_data_mask   ;
  input                                           std__pe8__lane24_strm1_data_valid  ;

  output                                          pe8__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane25_strm0_data_mask   ;
  input                                           std__pe8__lane25_strm0_data_valid  ;

  output                                          pe8__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane25_strm1_data_mask   ;
  input                                           std__pe8__lane25_strm1_data_valid  ;

  output                                          pe8__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane26_strm0_data_mask   ;
  input                                           std__pe8__lane26_strm0_data_valid  ;

  output                                          pe8__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane26_strm1_data_mask   ;
  input                                           std__pe8__lane26_strm1_data_valid  ;

  output                                          pe8__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane27_strm0_data_mask   ;
  input                                           std__pe8__lane27_strm0_data_valid  ;

  output                                          pe8__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane27_strm1_data_mask   ;
  input                                           std__pe8__lane27_strm1_data_valid  ;

  output                                          pe8__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane28_strm0_data_mask   ;
  input                                           std__pe8__lane28_strm0_data_valid  ;

  output                                          pe8__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane28_strm1_data_mask   ;
  input                                           std__pe8__lane28_strm1_data_valid  ;

  output                                          pe8__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane29_strm0_data_mask   ;
  input                                           std__pe8__lane29_strm0_data_valid  ;

  output                                          pe8__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane29_strm1_data_mask   ;
  input                                           std__pe8__lane29_strm1_data_valid  ;

  output                                          pe8__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane30_strm0_data_mask   ;
  input                                           std__pe8__lane30_strm0_data_valid  ;

  output                                          pe8__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane30_strm1_data_mask   ;
  input                                           std__pe8__lane30_strm1_data_valid  ;

  output                                          pe8__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane31_strm0_data_mask   ;
  input                                           std__pe8__lane31_strm0_data_valid  ;

  output                                          pe8__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe8__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe8__lane31_strm1_data_mask   ;
  input                                           std__pe8__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe9__peId                ;
  input                                         sys__pe9__allSynchronized     ;
  output                                        pe9__sys__thisSynchronized    ;
  output                                        pe9__sys__ready               ;
  output                                        pe9__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe9__oob_cntl            ;
  input                                         std__pe9__oob_valid           ;
  output                                        pe9__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe9__oob_type            ;
  output                                          pe9__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane0_strm0_data_mask   ;
  input                                           std__pe9__lane0_strm0_data_valid  ;

  output                                          pe9__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane0_strm1_data_mask   ;
  input                                           std__pe9__lane0_strm1_data_valid  ;

  output                                          pe9__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane1_strm0_data_mask   ;
  input                                           std__pe9__lane1_strm0_data_valid  ;

  output                                          pe9__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane1_strm1_data_mask   ;
  input                                           std__pe9__lane1_strm1_data_valid  ;

  output                                          pe9__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane2_strm0_data_mask   ;
  input                                           std__pe9__lane2_strm0_data_valid  ;

  output                                          pe9__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane2_strm1_data_mask   ;
  input                                           std__pe9__lane2_strm1_data_valid  ;

  output                                          pe9__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane3_strm0_data_mask   ;
  input                                           std__pe9__lane3_strm0_data_valid  ;

  output                                          pe9__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane3_strm1_data_mask   ;
  input                                           std__pe9__lane3_strm1_data_valid  ;

  output                                          pe9__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane4_strm0_data_mask   ;
  input                                           std__pe9__lane4_strm0_data_valid  ;

  output                                          pe9__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane4_strm1_data_mask   ;
  input                                           std__pe9__lane4_strm1_data_valid  ;

  output                                          pe9__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane5_strm0_data_mask   ;
  input                                           std__pe9__lane5_strm0_data_valid  ;

  output                                          pe9__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane5_strm1_data_mask   ;
  input                                           std__pe9__lane5_strm1_data_valid  ;

  output                                          pe9__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane6_strm0_data_mask   ;
  input                                           std__pe9__lane6_strm0_data_valid  ;

  output                                          pe9__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane6_strm1_data_mask   ;
  input                                           std__pe9__lane6_strm1_data_valid  ;

  output                                          pe9__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane7_strm0_data_mask   ;
  input                                           std__pe9__lane7_strm0_data_valid  ;

  output                                          pe9__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane7_strm1_data_mask   ;
  input                                           std__pe9__lane7_strm1_data_valid  ;

  output                                          pe9__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane8_strm0_data_mask   ;
  input                                           std__pe9__lane8_strm0_data_valid  ;

  output                                          pe9__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane8_strm1_data_mask   ;
  input                                           std__pe9__lane8_strm1_data_valid  ;

  output                                          pe9__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane9_strm0_data_mask   ;
  input                                           std__pe9__lane9_strm0_data_valid  ;

  output                                          pe9__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane9_strm1_data_mask   ;
  input                                           std__pe9__lane9_strm1_data_valid  ;

  output                                          pe9__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane10_strm0_data_mask   ;
  input                                           std__pe9__lane10_strm0_data_valid  ;

  output                                          pe9__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane10_strm1_data_mask   ;
  input                                           std__pe9__lane10_strm1_data_valid  ;

  output                                          pe9__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane11_strm0_data_mask   ;
  input                                           std__pe9__lane11_strm0_data_valid  ;

  output                                          pe9__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane11_strm1_data_mask   ;
  input                                           std__pe9__lane11_strm1_data_valid  ;

  output                                          pe9__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane12_strm0_data_mask   ;
  input                                           std__pe9__lane12_strm0_data_valid  ;

  output                                          pe9__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane12_strm1_data_mask   ;
  input                                           std__pe9__lane12_strm1_data_valid  ;

  output                                          pe9__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane13_strm0_data_mask   ;
  input                                           std__pe9__lane13_strm0_data_valid  ;

  output                                          pe9__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane13_strm1_data_mask   ;
  input                                           std__pe9__lane13_strm1_data_valid  ;

  output                                          pe9__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane14_strm0_data_mask   ;
  input                                           std__pe9__lane14_strm0_data_valid  ;

  output                                          pe9__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane14_strm1_data_mask   ;
  input                                           std__pe9__lane14_strm1_data_valid  ;

  output                                          pe9__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane15_strm0_data_mask   ;
  input                                           std__pe9__lane15_strm0_data_valid  ;

  output                                          pe9__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane15_strm1_data_mask   ;
  input                                           std__pe9__lane15_strm1_data_valid  ;

  output                                          pe9__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane16_strm0_data_mask   ;
  input                                           std__pe9__lane16_strm0_data_valid  ;

  output                                          pe9__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane16_strm1_data_mask   ;
  input                                           std__pe9__lane16_strm1_data_valid  ;

  output                                          pe9__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane17_strm0_data_mask   ;
  input                                           std__pe9__lane17_strm0_data_valid  ;

  output                                          pe9__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane17_strm1_data_mask   ;
  input                                           std__pe9__lane17_strm1_data_valid  ;

  output                                          pe9__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane18_strm0_data_mask   ;
  input                                           std__pe9__lane18_strm0_data_valid  ;

  output                                          pe9__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane18_strm1_data_mask   ;
  input                                           std__pe9__lane18_strm1_data_valid  ;

  output                                          pe9__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane19_strm0_data_mask   ;
  input                                           std__pe9__lane19_strm0_data_valid  ;

  output                                          pe9__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane19_strm1_data_mask   ;
  input                                           std__pe9__lane19_strm1_data_valid  ;

  output                                          pe9__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane20_strm0_data_mask   ;
  input                                           std__pe9__lane20_strm0_data_valid  ;

  output                                          pe9__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane20_strm1_data_mask   ;
  input                                           std__pe9__lane20_strm1_data_valid  ;

  output                                          pe9__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane21_strm0_data_mask   ;
  input                                           std__pe9__lane21_strm0_data_valid  ;

  output                                          pe9__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane21_strm1_data_mask   ;
  input                                           std__pe9__lane21_strm1_data_valid  ;

  output                                          pe9__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane22_strm0_data_mask   ;
  input                                           std__pe9__lane22_strm0_data_valid  ;

  output                                          pe9__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane22_strm1_data_mask   ;
  input                                           std__pe9__lane22_strm1_data_valid  ;

  output                                          pe9__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane23_strm0_data_mask   ;
  input                                           std__pe9__lane23_strm0_data_valid  ;

  output                                          pe9__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane23_strm1_data_mask   ;
  input                                           std__pe9__lane23_strm1_data_valid  ;

  output                                          pe9__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane24_strm0_data_mask   ;
  input                                           std__pe9__lane24_strm0_data_valid  ;

  output                                          pe9__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane24_strm1_data_mask   ;
  input                                           std__pe9__lane24_strm1_data_valid  ;

  output                                          pe9__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane25_strm0_data_mask   ;
  input                                           std__pe9__lane25_strm0_data_valid  ;

  output                                          pe9__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane25_strm1_data_mask   ;
  input                                           std__pe9__lane25_strm1_data_valid  ;

  output                                          pe9__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane26_strm0_data_mask   ;
  input                                           std__pe9__lane26_strm0_data_valid  ;

  output                                          pe9__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane26_strm1_data_mask   ;
  input                                           std__pe9__lane26_strm1_data_valid  ;

  output                                          pe9__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane27_strm0_data_mask   ;
  input                                           std__pe9__lane27_strm0_data_valid  ;

  output                                          pe9__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane27_strm1_data_mask   ;
  input                                           std__pe9__lane27_strm1_data_valid  ;

  output                                          pe9__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane28_strm0_data_mask   ;
  input                                           std__pe9__lane28_strm0_data_valid  ;

  output                                          pe9__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane28_strm1_data_mask   ;
  input                                           std__pe9__lane28_strm1_data_valid  ;

  output                                          pe9__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane29_strm0_data_mask   ;
  input                                           std__pe9__lane29_strm0_data_valid  ;

  output                                          pe9__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane29_strm1_data_mask   ;
  input                                           std__pe9__lane29_strm1_data_valid  ;

  output                                          pe9__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane30_strm0_data_mask   ;
  input                                           std__pe9__lane30_strm0_data_valid  ;

  output                                          pe9__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane30_strm1_data_mask   ;
  input                                           std__pe9__lane30_strm1_data_valid  ;

  output                                          pe9__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane31_strm0_data_mask   ;
  input                                           std__pe9__lane31_strm0_data_valid  ;

  output                                          pe9__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe9__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe9__lane31_strm1_data_mask   ;
  input                                           std__pe9__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe10__peId                ;
  input                                         sys__pe10__allSynchronized     ;
  output                                        pe10__sys__thisSynchronized    ;
  output                                        pe10__sys__ready               ;
  output                                        pe10__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe10__oob_cntl            ;
  input                                         std__pe10__oob_valid           ;
  output                                        pe10__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe10__oob_type            ;
  output                                          pe10__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane0_strm0_data_mask   ;
  input                                           std__pe10__lane0_strm0_data_valid  ;

  output                                          pe10__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane0_strm1_data_mask   ;
  input                                           std__pe10__lane0_strm1_data_valid  ;

  output                                          pe10__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane1_strm0_data_mask   ;
  input                                           std__pe10__lane1_strm0_data_valid  ;

  output                                          pe10__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane1_strm1_data_mask   ;
  input                                           std__pe10__lane1_strm1_data_valid  ;

  output                                          pe10__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane2_strm0_data_mask   ;
  input                                           std__pe10__lane2_strm0_data_valid  ;

  output                                          pe10__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane2_strm1_data_mask   ;
  input                                           std__pe10__lane2_strm1_data_valid  ;

  output                                          pe10__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane3_strm0_data_mask   ;
  input                                           std__pe10__lane3_strm0_data_valid  ;

  output                                          pe10__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane3_strm1_data_mask   ;
  input                                           std__pe10__lane3_strm1_data_valid  ;

  output                                          pe10__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane4_strm0_data_mask   ;
  input                                           std__pe10__lane4_strm0_data_valid  ;

  output                                          pe10__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane4_strm1_data_mask   ;
  input                                           std__pe10__lane4_strm1_data_valid  ;

  output                                          pe10__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane5_strm0_data_mask   ;
  input                                           std__pe10__lane5_strm0_data_valid  ;

  output                                          pe10__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane5_strm1_data_mask   ;
  input                                           std__pe10__lane5_strm1_data_valid  ;

  output                                          pe10__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane6_strm0_data_mask   ;
  input                                           std__pe10__lane6_strm0_data_valid  ;

  output                                          pe10__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane6_strm1_data_mask   ;
  input                                           std__pe10__lane6_strm1_data_valid  ;

  output                                          pe10__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane7_strm0_data_mask   ;
  input                                           std__pe10__lane7_strm0_data_valid  ;

  output                                          pe10__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane7_strm1_data_mask   ;
  input                                           std__pe10__lane7_strm1_data_valid  ;

  output                                          pe10__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane8_strm0_data_mask   ;
  input                                           std__pe10__lane8_strm0_data_valid  ;

  output                                          pe10__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane8_strm1_data_mask   ;
  input                                           std__pe10__lane8_strm1_data_valid  ;

  output                                          pe10__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane9_strm0_data_mask   ;
  input                                           std__pe10__lane9_strm0_data_valid  ;

  output                                          pe10__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane9_strm1_data_mask   ;
  input                                           std__pe10__lane9_strm1_data_valid  ;

  output                                          pe10__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane10_strm0_data_mask   ;
  input                                           std__pe10__lane10_strm0_data_valid  ;

  output                                          pe10__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane10_strm1_data_mask   ;
  input                                           std__pe10__lane10_strm1_data_valid  ;

  output                                          pe10__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane11_strm0_data_mask   ;
  input                                           std__pe10__lane11_strm0_data_valid  ;

  output                                          pe10__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane11_strm1_data_mask   ;
  input                                           std__pe10__lane11_strm1_data_valid  ;

  output                                          pe10__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane12_strm0_data_mask   ;
  input                                           std__pe10__lane12_strm0_data_valid  ;

  output                                          pe10__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane12_strm1_data_mask   ;
  input                                           std__pe10__lane12_strm1_data_valid  ;

  output                                          pe10__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane13_strm0_data_mask   ;
  input                                           std__pe10__lane13_strm0_data_valid  ;

  output                                          pe10__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane13_strm1_data_mask   ;
  input                                           std__pe10__lane13_strm1_data_valid  ;

  output                                          pe10__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane14_strm0_data_mask   ;
  input                                           std__pe10__lane14_strm0_data_valid  ;

  output                                          pe10__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane14_strm1_data_mask   ;
  input                                           std__pe10__lane14_strm1_data_valid  ;

  output                                          pe10__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane15_strm0_data_mask   ;
  input                                           std__pe10__lane15_strm0_data_valid  ;

  output                                          pe10__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane15_strm1_data_mask   ;
  input                                           std__pe10__lane15_strm1_data_valid  ;

  output                                          pe10__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane16_strm0_data_mask   ;
  input                                           std__pe10__lane16_strm0_data_valid  ;

  output                                          pe10__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane16_strm1_data_mask   ;
  input                                           std__pe10__lane16_strm1_data_valid  ;

  output                                          pe10__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane17_strm0_data_mask   ;
  input                                           std__pe10__lane17_strm0_data_valid  ;

  output                                          pe10__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane17_strm1_data_mask   ;
  input                                           std__pe10__lane17_strm1_data_valid  ;

  output                                          pe10__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane18_strm0_data_mask   ;
  input                                           std__pe10__lane18_strm0_data_valid  ;

  output                                          pe10__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane18_strm1_data_mask   ;
  input                                           std__pe10__lane18_strm1_data_valid  ;

  output                                          pe10__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane19_strm0_data_mask   ;
  input                                           std__pe10__lane19_strm0_data_valid  ;

  output                                          pe10__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane19_strm1_data_mask   ;
  input                                           std__pe10__lane19_strm1_data_valid  ;

  output                                          pe10__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane20_strm0_data_mask   ;
  input                                           std__pe10__lane20_strm0_data_valid  ;

  output                                          pe10__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane20_strm1_data_mask   ;
  input                                           std__pe10__lane20_strm1_data_valid  ;

  output                                          pe10__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane21_strm0_data_mask   ;
  input                                           std__pe10__lane21_strm0_data_valid  ;

  output                                          pe10__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane21_strm1_data_mask   ;
  input                                           std__pe10__lane21_strm1_data_valid  ;

  output                                          pe10__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane22_strm0_data_mask   ;
  input                                           std__pe10__lane22_strm0_data_valid  ;

  output                                          pe10__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane22_strm1_data_mask   ;
  input                                           std__pe10__lane22_strm1_data_valid  ;

  output                                          pe10__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane23_strm0_data_mask   ;
  input                                           std__pe10__lane23_strm0_data_valid  ;

  output                                          pe10__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane23_strm1_data_mask   ;
  input                                           std__pe10__lane23_strm1_data_valid  ;

  output                                          pe10__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane24_strm0_data_mask   ;
  input                                           std__pe10__lane24_strm0_data_valid  ;

  output                                          pe10__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane24_strm1_data_mask   ;
  input                                           std__pe10__lane24_strm1_data_valid  ;

  output                                          pe10__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane25_strm0_data_mask   ;
  input                                           std__pe10__lane25_strm0_data_valid  ;

  output                                          pe10__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane25_strm1_data_mask   ;
  input                                           std__pe10__lane25_strm1_data_valid  ;

  output                                          pe10__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane26_strm0_data_mask   ;
  input                                           std__pe10__lane26_strm0_data_valid  ;

  output                                          pe10__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane26_strm1_data_mask   ;
  input                                           std__pe10__lane26_strm1_data_valid  ;

  output                                          pe10__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane27_strm0_data_mask   ;
  input                                           std__pe10__lane27_strm0_data_valid  ;

  output                                          pe10__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane27_strm1_data_mask   ;
  input                                           std__pe10__lane27_strm1_data_valid  ;

  output                                          pe10__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane28_strm0_data_mask   ;
  input                                           std__pe10__lane28_strm0_data_valid  ;

  output                                          pe10__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane28_strm1_data_mask   ;
  input                                           std__pe10__lane28_strm1_data_valid  ;

  output                                          pe10__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane29_strm0_data_mask   ;
  input                                           std__pe10__lane29_strm0_data_valid  ;

  output                                          pe10__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane29_strm1_data_mask   ;
  input                                           std__pe10__lane29_strm1_data_valid  ;

  output                                          pe10__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane30_strm0_data_mask   ;
  input                                           std__pe10__lane30_strm0_data_valid  ;

  output                                          pe10__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane30_strm1_data_mask   ;
  input                                           std__pe10__lane30_strm1_data_valid  ;

  output                                          pe10__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane31_strm0_data_mask   ;
  input                                           std__pe10__lane31_strm0_data_valid  ;

  output                                          pe10__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe10__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe10__lane31_strm1_data_mask   ;
  input                                           std__pe10__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe11__peId                ;
  input                                         sys__pe11__allSynchronized     ;
  output                                        pe11__sys__thisSynchronized    ;
  output                                        pe11__sys__ready               ;
  output                                        pe11__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe11__oob_cntl            ;
  input                                         std__pe11__oob_valid           ;
  output                                        pe11__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe11__oob_type            ;
  output                                          pe11__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane0_strm0_data_mask   ;
  input                                           std__pe11__lane0_strm0_data_valid  ;

  output                                          pe11__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane0_strm1_data_mask   ;
  input                                           std__pe11__lane0_strm1_data_valid  ;

  output                                          pe11__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane1_strm0_data_mask   ;
  input                                           std__pe11__lane1_strm0_data_valid  ;

  output                                          pe11__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane1_strm1_data_mask   ;
  input                                           std__pe11__lane1_strm1_data_valid  ;

  output                                          pe11__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane2_strm0_data_mask   ;
  input                                           std__pe11__lane2_strm0_data_valid  ;

  output                                          pe11__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane2_strm1_data_mask   ;
  input                                           std__pe11__lane2_strm1_data_valid  ;

  output                                          pe11__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane3_strm0_data_mask   ;
  input                                           std__pe11__lane3_strm0_data_valid  ;

  output                                          pe11__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane3_strm1_data_mask   ;
  input                                           std__pe11__lane3_strm1_data_valid  ;

  output                                          pe11__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane4_strm0_data_mask   ;
  input                                           std__pe11__lane4_strm0_data_valid  ;

  output                                          pe11__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane4_strm1_data_mask   ;
  input                                           std__pe11__lane4_strm1_data_valid  ;

  output                                          pe11__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane5_strm0_data_mask   ;
  input                                           std__pe11__lane5_strm0_data_valid  ;

  output                                          pe11__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane5_strm1_data_mask   ;
  input                                           std__pe11__lane5_strm1_data_valid  ;

  output                                          pe11__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane6_strm0_data_mask   ;
  input                                           std__pe11__lane6_strm0_data_valid  ;

  output                                          pe11__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane6_strm1_data_mask   ;
  input                                           std__pe11__lane6_strm1_data_valid  ;

  output                                          pe11__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane7_strm0_data_mask   ;
  input                                           std__pe11__lane7_strm0_data_valid  ;

  output                                          pe11__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane7_strm1_data_mask   ;
  input                                           std__pe11__lane7_strm1_data_valid  ;

  output                                          pe11__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane8_strm0_data_mask   ;
  input                                           std__pe11__lane8_strm0_data_valid  ;

  output                                          pe11__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane8_strm1_data_mask   ;
  input                                           std__pe11__lane8_strm1_data_valid  ;

  output                                          pe11__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane9_strm0_data_mask   ;
  input                                           std__pe11__lane9_strm0_data_valid  ;

  output                                          pe11__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane9_strm1_data_mask   ;
  input                                           std__pe11__lane9_strm1_data_valid  ;

  output                                          pe11__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane10_strm0_data_mask   ;
  input                                           std__pe11__lane10_strm0_data_valid  ;

  output                                          pe11__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane10_strm1_data_mask   ;
  input                                           std__pe11__lane10_strm1_data_valid  ;

  output                                          pe11__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane11_strm0_data_mask   ;
  input                                           std__pe11__lane11_strm0_data_valid  ;

  output                                          pe11__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane11_strm1_data_mask   ;
  input                                           std__pe11__lane11_strm1_data_valid  ;

  output                                          pe11__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane12_strm0_data_mask   ;
  input                                           std__pe11__lane12_strm0_data_valid  ;

  output                                          pe11__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane12_strm1_data_mask   ;
  input                                           std__pe11__lane12_strm1_data_valid  ;

  output                                          pe11__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane13_strm0_data_mask   ;
  input                                           std__pe11__lane13_strm0_data_valid  ;

  output                                          pe11__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane13_strm1_data_mask   ;
  input                                           std__pe11__lane13_strm1_data_valid  ;

  output                                          pe11__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane14_strm0_data_mask   ;
  input                                           std__pe11__lane14_strm0_data_valid  ;

  output                                          pe11__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane14_strm1_data_mask   ;
  input                                           std__pe11__lane14_strm1_data_valid  ;

  output                                          pe11__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane15_strm0_data_mask   ;
  input                                           std__pe11__lane15_strm0_data_valid  ;

  output                                          pe11__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane15_strm1_data_mask   ;
  input                                           std__pe11__lane15_strm1_data_valid  ;

  output                                          pe11__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane16_strm0_data_mask   ;
  input                                           std__pe11__lane16_strm0_data_valid  ;

  output                                          pe11__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane16_strm1_data_mask   ;
  input                                           std__pe11__lane16_strm1_data_valid  ;

  output                                          pe11__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane17_strm0_data_mask   ;
  input                                           std__pe11__lane17_strm0_data_valid  ;

  output                                          pe11__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane17_strm1_data_mask   ;
  input                                           std__pe11__lane17_strm1_data_valid  ;

  output                                          pe11__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane18_strm0_data_mask   ;
  input                                           std__pe11__lane18_strm0_data_valid  ;

  output                                          pe11__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane18_strm1_data_mask   ;
  input                                           std__pe11__lane18_strm1_data_valid  ;

  output                                          pe11__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane19_strm0_data_mask   ;
  input                                           std__pe11__lane19_strm0_data_valid  ;

  output                                          pe11__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane19_strm1_data_mask   ;
  input                                           std__pe11__lane19_strm1_data_valid  ;

  output                                          pe11__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane20_strm0_data_mask   ;
  input                                           std__pe11__lane20_strm0_data_valid  ;

  output                                          pe11__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane20_strm1_data_mask   ;
  input                                           std__pe11__lane20_strm1_data_valid  ;

  output                                          pe11__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane21_strm0_data_mask   ;
  input                                           std__pe11__lane21_strm0_data_valid  ;

  output                                          pe11__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane21_strm1_data_mask   ;
  input                                           std__pe11__lane21_strm1_data_valid  ;

  output                                          pe11__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane22_strm0_data_mask   ;
  input                                           std__pe11__lane22_strm0_data_valid  ;

  output                                          pe11__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane22_strm1_data_mask   ;
  input                                           std__pe11__lane22_strm1_data_valid  ;

  output                                          pe11__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane23_strm0_data_mask   ;
  input                                           std__pe11__lane23_strm0_data_valid  ;

  output                                          pe11__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane23_strm1_data_mask   ;
  input                                           std__pe11__lane23_strm1_data_valid  ;

  output                                          pe11__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane24_strm0_data_mask   ;
  input                                           std__pe11__lane24_strm0_data_valid  ;

  output                                          pe11__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane24_strm1_data_mask   ;
  input                                           std__pe11__lane24_strm1_data_valid  ;

  output                                          pe11__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane25_strm0_data_mask   ;
  input                                           std__pe11__lane25_strm0_data_valid  ;

  output                                          pe11__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane25_strm1_data_mask   ;
  input                                           std__pe11__lane25_strm1_data_valid  ;

  output                                          pe11__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane26_strm0_data_mask   ;
  input                                           std__pe11__lane26_strm0_data_valid  ;

  output                                          pe11__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane26_strm1_data_mask   ;
  input                                           std__pe11__lane26_strm1_data_valid  ;

  output                                          pe11__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane27_strm0_data_mask   ;
  input                                           std__pe11__lane27_strm0_data_valid  ;

  output                                          pe11__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane27_strm1_data_mask   ;
  input                                           std__pe11__lane27_strm1_data_valid  ;

  output                                          pe11__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane28_strm0_data_mask   ;
  input                                           std__pe11__lane28_strm0_data_valid  ;

  output                                          pe11__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane28_strm1_data_mask   ;
  input                                           std__pe11__lane28_strm1_data_valid  ;

  output                                          pe11__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane29_strm0_data_mask   ;
  input                                           std__pe11__lane29_strm0_data_valid  ;

  output                                          pe11__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane29_strm1_data_mask   ;
  input                                           std__pe11__lane29_strm1_data_valid  ;

  output                                          pe11__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane30_strm0_data_mask   ;
  input                                           std__pe11__lane30_strm0_data_valid  ;

  output                                          pe11__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane30_strm1_data_mask   ;
  input                                           std__pe11__lane30_strm1_data_valid  ;

  output                                          pe11__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane31_strm0_data_mask   ;
  input                                           std__pe11__lane31_strm0_data_valid  ;

  output                                          pe11__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe11__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe11__lane31_strm1_data_mask   ;
  input                                           std__pe11__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe12__peId                ;
  input                                         sys__pe12__allSynchronized     ;
  output                                        pe12__sys__thisSynchronized    ;
  output                                        pe12__sys__ready               ;
  output                                        pe12__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe12__oob_cntl            ;
  input                                         std__pe12__oob_valid           ;
  output                                        pe12__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe12__oob_type            ;
  output                                          pe12__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane0_strm0_data_mask   ;
  input                                           std__pe12__lane0_strm0_data_valid  ;

  output                                          pe12__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane0_strm1_data_mask   ;
  input                                           std__pe12__lane0_strm1_data_valid  ;

  output                                          pe12__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane1_strm0_data_mask   ;
  input                                           std__pe12__lane1_strm0_data_valid  ;

  output                                          pe12__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane1_strm1_data_mask   ;
  input                                           std__pe12__lane1_strm1_data_valid  ;

  output                                          pe12__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane2_strm0_data_mask   ;
  input                                           std__pe12__lane2_strm0_data_valid  ;

  output                                          pe12__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane2_strm1_data_mask   ;
  input                                           std__pe12__lane2_strm1_data_valid  ;

  output                                          pe12__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane3_strm0_data_mask   ;
  input                                           std__pe12__lane3_strm0_data_valid  ;

  output                                          pe12__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane3_strm1_data_mask   ;
  input                                           std__pe12__lane3_strm1_data_valid  ;

  output                                          pe12__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane4_strm0_data_mask   ;
  input                                           std__pe12__lane4_strm0_data_valid  ;

  output                                          pe12__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane4_strm1_data_mask   ;
  input                                           std__pe12__lane4_strm1_data_valid  ;

  output                                          pe12__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane5_strm0_data_mask   ;
  input                                           std__pe12__lane5_strm0_data_valid  ;

  output                                          pe12__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane5_strm1_data_mask   ;
  input                                           std__pe12__lane5_strm1_data_valid  ;

  output                                          pe12__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane6_strm0_data_mask   ;
  input                                           std__pe12__lane6_strm0_data_valid  ;

  output                                          pe12__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane6_strm1_data_mask   ;
  input                                           std__pe12__lane6_strm1_data_valid  ;

  output                                          pe12__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane7_strm0_data_mask   ;
  input                                           std__pe12__lane7_strm0_data_valid  ;

  output                                          pe12__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane7_strm1_data_mask   ;
  input                                           std__pe12__lane7_strm1_data_valid  ;

  output                                          pe12__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane8_strm0_data_mask   ;
  input                                           std__pe12__lane8_strm0_data_valid  ;

  output                                          pe12__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane8_strm1_data_mask   ;
  input                                           std__pe12__lane8_strm1_data_valid  ;

  output                                          pe12__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane9_strm0_data_mask   ;
  input                                           std__pe12__lane9_strm0_data_valid  ;

  output                                          pe12__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane9_strm1_data_mask   ;
  input                                           std__pe12__lane9_strm1_data_valid  ;

  output                                          pe12__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane10_strm0_data_mask   ;
  input                                           std__pe12__lane10_strm0_data_valid  ;

  output                                          pe12__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane10_strm1_data_mask   ;
  input                                           std__pe12__lane10_strm1_data_valid  ;

  output                                          pe12__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane11_strm0_data_mask   ;
  input                                           std__pe12__lane11_strm0_data_valid  ;

  output                                          pe12__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane11_strm1_data_mask   ;
  input                                           std__pe12__lane11_strm1_data_valid  ;

  output                                          pe12__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane12_strm0_data_mask   ;
  input                                           std__pe12__lane12_strm0_data_valid  ;

  output                                          pe12__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane12_strm1_data_mask   ;
  input                                           std__pe12__lane12_strm1_data_valid  ;

  output                                          pe12__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane13_strm0_data_mask   ;
  input                                           std__pe12__lane13_strm0_data_valid  ;

  output                                          pe12__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane13_strm1_data_mask   ;
  input                                           std__pe12__lane13_strm1_data_valid  ;

  output                                          pe12__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane14_strm0_data_mask   ;
  input                                           std__pe12__lane14_strm0_data_valid  ;

  output                                          pe12__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane14_strm1_data_mask   ;
  input                                           std__pe12__lane14_strm1_data_valid  ;

  output                                          pe12__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane15_strm0_data_mask   ;
  input                                           std__pe12__lane15_strm0_data_valid  ;

  output                                          pe12__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane15_strm1_data_mask   ;
  input                                           std__pe12__lane15_strm1_data_valid  ;

  output                                          pe12__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane16_strm0_data_mask   ;
  input                                           std__pe12__lane16_strm0_data_valid  ;

  output                                          pe12__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane16_strm1_data_mask   ;
  input                                           std__pe12__lane16_strm1_data_valid  ;

  output                                          pe12__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane17_strm0_data_mask   ;
  input                                           std__pe12__lane17_strm0_data_valid  ;

  output                                          pe12__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane17_strm1_data_mask   ;
  input                                           std__pe12__lane17_strm1_data_valid  ;

  output                                          pe12__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane18_strm0_data_mask   ;
  input                                           std__pe12__lane18_strm0_data_valid  ;

  output                                          pe12__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane18_strm1_data_mask   ;
  input                                           std__pe12__lane18_strm1_data_valid  ;

  output                                          pe12__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane19_strm0_data_mask   ;
  input                                           std__pe12__lane19_strm0_data_valid  ;

  output                                          pe12__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane19_strm1_data_mask   ;
  input                                           std__pe12__lane19_strm1_data_valid  ;

  output                                          pe12__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane20_strm0_data_mask   ;
  input                                           std__pe12__lane20_strm0_data_valid  ;

  output                                          pe12__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane20_strm1_data_mask   ;
  input                                           std__pe12__lane20_strm1_data_valid  ;

  output                                          pe12__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane21_strm0_data_mask   ;
  input                                           std__pe12__lane21_strm0_data_valid  ;

  output                                          pe12__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane21_strm1_data_mask   ;
  input                                           std__pe12__lane21_strm1_data_valid  ;

  output                                          pe12__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane22_strm0_data_mask   ;
  input                                           std__pe12__lane22_strm0_data_valid  ;

  output                                          pe12__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane22_strm1_data_mask   ;
  input                                           std__pe12__lane22_strm1_data_valid  ;

  output                                          pe12__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane23_strm0_data_mask   ;
  input                                           std__pe12__lane23_strm0_data_valid  ;

  output                                          pe12__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane23_strm1_data_mask   ;
  input                                           std__pe12__lane23_strm1_data_valid  ;

  output                                          pe12__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane24_strm0_data_mask   ;
  input                                           std__pe12__lane24_strm0_data_valid  ;

  output                                          pe12__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane24_strm1_data_mask   ;
  input                                           std__pe12__lane24_strm1_data_valid  ;

  output                                          pe12__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane25_strm0_data_mask   ;
  input                                           std__pe12__lane25_strm0_data_valid  ;

  output                                          pe12__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane25_strm1_data_mask   ;
  input                                           std__pe12__lane25_strm1_data_valid  ;

  output                                          pe12__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane26_strm0_data_mask   ;
  input                                           std__pe12__lane26_strm0_data_valid  ;

  output                                          pe12__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane26_strm1_data_mask   ;
  input                                           std__pe12__lane26_strm1_data_valid  ;

  output                                          pe12__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane27_strm0_data_mask   ;
  input                                           std__pe12__lane27_strm0_data_valid  ;

  output                                          pe12__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane27_strm1_data_mask   ;
  input                                           std__pe12__lane27_strm1_data_valid  ;

  output                                          pe12__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane28_strm0_data_mask   ;
  input                                           std__pe12__lane28_strm0_data_valid  ;

  output                                          pe12__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane28_strm1_data_mask   ;
  input                                           std__pe12__lane28_strm1_data_valid  ;

  output                                          pe12__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane29_strm0_data_mask   ;
  input                                           std__pe12__lane29_strm0_data_valid  ;

  output                                          pe12__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane29_strm1_data_mask   ;
  input                                           std__pe12__lane29_strm1_data_valid  ;

  output                                          pe12__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane30_strm0_data_mask   ;
  input                                           std__pe12__lane30_strm0_data_valid  ;

  output                                          pe12__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane30_strm1_data_mask   ;
  input                                           std__pe12__lane30_strm1_data_valid  ;

  output                                          pe12__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane31_strm0_data_mask   ;
  input                                           std__pe12__lane31_strm0_data_valid  ;

  output                                          pe12__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe12__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe12__lane31_strm1_data_mask   ;
  input                                           std__pe12__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe13__peId                ;
  input                                         sys__pe13__allSynchronized     ;
  output                                        pe13__sys__thisSynchronized    ;
  output                                        pe13__sys__ready               ;
  output                                        pe13__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe13__oob_cntl            ;
  input                                         std__pe13__oob_valid           ;
  output                                        pe13__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe13__oob_type            ;
  output                                          pe13__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane0_strm0_data_mask   ;
  input                                           std__pe13__lane0_strm0_data_valid  ;

  output                                          pe13__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane0_strm1_data_mask   ;
  input                                           std__pe13__lane0_strm1_data_valid  ;

  output                                          pe13__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane1_strm0_data_mask   ;
  input                                           std__pe13__lane1_strm0_data_valid  ;

  output                                          pe13__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane1_strm1_data_mask   ;
  input                                           std__pe13__lane1_strm1_data_valid  ;

  output                                          pe13__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane2_strm0_data_mask   ;
  input                                           std__pe13__lane2_strm0_data_valid  ;

  output                                          pe13__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane2_strm1_data_mask   ;
  input                                           std__pe13__lane2_strm1_data_valid  ;

  output                                          pe13__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane3_strm0_data_mask   ;
  input                                           std__pe13__lane3_strm0_data_valid  ;

  output                                          pe13__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane3_strm1_data_mask   ;
  input                                           std__pe13__lane3_strm1_data_valid  ;

  output                                          pe13__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane4_strm0_data_mask   ;
  input                                           std__pe13__lane4_strm0_data_valid  ;

  output                                          pe13__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane4_strm1_data_mask   ;
  input                                           std__pe13__lane4_strm1_data_valid  ;

  output                                          pe13__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane5_strm0_data_mask   ;
  input                                           std__pe13__lane5_strm0_data_valid  ;

  output                                          pe13__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane5_strm1_data_mask   ;
  input                                           std__pe13__lane5_strm1_data_valid  ;

  output                                          pe13__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane6_strm0_data_mask   ;
  input                                           std__pe13__lane6_strm0_data_valid  ;

  output                                          pe13__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane6_strm1_data_mask   ;
  input                                           std__pe13__lane6_strm1_data_valid  ;

  output                                          pe13__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane7_strm0_data_mask   ;
  input                                           std__pe13__lane7_strm0_data_valid  ;

  output                                          pe13__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane7_strm1_data_mask   ;
  input                                           std__pe13__lane7_strm1_data_valid  ;

  output                                          pe13__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane8_strm0_data_mask   ;
  input                                           std__pe13__lane8_strm0_data_valid  ;

  output                                          pe13__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane8_strm1_data_mask   ;
  input                                           std__pe13__lane8_strm1_data_valid  ;

  output                                          pe13__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane9_strm0_data_mask   ;
  input                                           std__pe13__lane9_strm0_data_valid  ;

  output                                          pe13__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane9_strm1_data_mask   ;
  input                                           std__pe13__lane9_strm1_data_valid  ;

  output                                          pe13__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane10_strm0_data_mask   ;
  input                                           std__pe13__lane10_strm0_data_valid  ;

  output                                          pe13__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane10_strm1_data_mask   ;
  input                                           std__pe13__lane10_strm1_data_valid  ;

  output                                          pe13__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane11_strm0_data_mask   ;
  input                                           std__pe13__lane11_strm0_data_valid  ;

  output                                          pe13__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane11_strm1_data_mask   ;
  input                                           std__pe13__lane11_strm1_data_valid  ;

  output                                          pe13__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane12_strm0_data_mask   ;
  input                                           std__pe13__lane12_strm0_data_valid  ;

  output                                          pe13__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane12_strm1_data_mask   ;
  input                                           std__pe13__lane12_strm1_data_valid  ;

  output                                          pe13__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane13_strm0_data_mask   ;
  input                                           std__pe13__lane13_strm0_data_valid  ;

  output                                          pe13__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane13_strm1_data_mask   ;
  input                                           std__pe13__lane13_strm1_data_valid  ;

  output                                          pe13__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane14_strm0_data_mask   ;
  input                                           std__pe13__lane14_strm0_data_valid  ;

  output                                          pe13__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane14_strm1_data_mask   ;
  input                                           std__pe13__lane14_strm1_data_valid  ;

  output                                          pe13__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane15_strm0_data_mask   ;
  input                                           std__pe13__lane15_strm0_data_valid  ;

  output                                          pe13__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane15_strm1_data_mask   ;
  input                                           std__pe13__lane15_strm1_data_valid  ;

  output                                          pe13__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane16_strm0_data_mask   ;
  input                                           std__pe13__lane16_strm0_data_valid  ;

  output                                          pe13__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane16_strm1_data_mask   ;
  input                                           std__pe13__lane16_strm1_data_valid  ;

  output                                          pe13__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane17_strm0_data_mask   ;
  input                                           std__pe13__lane17_strm0_data_valid  ;

  output                                          pe13__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane17_strm1_data_mask   ;
  input                                           std__pe13__lane17_strm1_data_valid  ;

  output                                          pe13__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane18_strm0_data_mask   ;
  input                                           std__pe13__lane18_strm0_data_valid  ;

  output                                          pe13__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane18_strm1_data_mask   ;
  input                                           std__pe13__lane18_strm1_data_valid  ;

  output                                          pe13__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane19_strm0_data_mask   ;
  input                                           std__pe13__lane19_strm0_data_valid  ;

  output                                          pe13__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane19_strm1_data_mask   ;
  input                                           std__pe13__lane19_strm1_data_valid  ;

  output                                          pe13__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane20_strm0_data_mask   ;
  input                                           std__pe13__lane20_strm0_data_valid  ;

  output                                          pe13__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane20_strm1_data_mask   ;
  input                                           std__pe13__lane20_strm1_data_valid  ;

  output                                          pe13__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane21_strm0_data_mask   ;
  input                                           std__pe13__lane21_strm0_data_valid  ;

  output                                          pe13__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane21_strm1_data_mask   ;
  input                                           std__pe13__lane21_strm1_data_valid  ;

  output                                          pe13__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane22_strm0_data_mask   ;
  input                                           std__pe13__lane22_strm0_data_valid  ;

  output                                          pe13__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane22_strm1_data_mask   ;
  input                                           std__pe13__lane22_strm1_data_valid  ;

  output                                          pe13__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane23_strm0_data_mask   ;
  input                                           std__pe13__lane23_strm0_data_valid  ;

  output                                          pe13__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane23_strm1_data_mask   ;
  input                                           std__pe13__lane23_strm1_data_valid  ;

  output                                          pe13__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane24_strm0_data_mask   ;
  input                                           std__pe13__lane24_strm0_data_valid  ;

  output                                          pe13__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane24_strm1_data_mask   ;
  input                                           std__pe13__lane24_strm1_data_valid  ;

  output                                          pe13__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane25_strm0_data_mask   ;
  input                                           std__pe13__lane25_strm0_data_valid  ;

  output                                          pe13__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane25_strm1_data_mask   ;
  input                                           std__pe13__lane25_strm1_data_valid  ;

  output                                          pe13__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane26_strm0_data_mask   ;
  input                                           std__pe13__lane26_strm0_data_valid  ;

  output                                          pe13__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane26_strm1_data_mask   ;
  input                                           std__pe13__lane26_strm1_data_valid  ;

  output                                          pe13__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane27_strm0_data_mask   ;
  input                                           std__pe13__lane27_strm0_data_valid  ;

  output                                          pe13__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane27_strm1_data_mask   ;
  input                                           std__pe13__lane27_strm1_data_valid  ;

  output                                          pe13__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane28_strm0_data_mask   ;
  input                                           std__pe13__lane28_strm0_data_valid  ;

  output                                          pe13__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane28_strm1_data_mask   ;
  input                                           std__pe13__lane28_strm1_data_valid  ;

  output                                          pe13__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane29_strm0_data_mask   ;
  input                                           std__pe13__lane29_strm0_data_valid  ;

  output                                          pe13__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane29_strm1_data_mask   ;
  input                                           std__pe13__lane29_strm1_data_valid  ;

  output                                          pe13__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane30_strm0_data_mask   ;
  input                                           std__pe13__lane30_strm0_data_valid  ;

  output                                          pe13__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane30_strm1_data_mask   ;
  input                                           std__pe13__lane30_strm1_data_valid  ;

  output                                          pe13__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane31_strm0_data_mask   ;
  input                                           std__pe13__lane31_strm0_data_valid  ;

  output                                          pe13__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe13__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe13__lane31_strm1_data_mask   ;
  input                                           std__pe13__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe14__peId                ;
  input                                         sys__pe14__allSynchronized     ;
  output                                        pe14__sys__thisSynchronized    ;
  output                                        pe14__sys__ready               ;
  output                                        pe14__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe14__oob_cntl            ;
  input                                         std__pe14__oob_valid           ;
  output                                        pe14__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe14__oob_type            ;
  output                                          pe14__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane0_strm0_data_mask   ;
  input                                           std__pe14__lane0_strm0_data_valid  ;

  output                                          pe14__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane0_strm1_data_mask   ;
  input                                           std__pe14__lane0_strm1_data_valid  ;

  output                                          pe14__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane1_strm0_data_mask   ;
  input                                           std__pe14__lane1_strm0_data_valid  ;

  output                                          pe14__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane1_strm1_data_mask   ;
  input                                           std__pe14__lane1_strm1_data_valid  ;

  output                                          pe14__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane2_strm0_data_mask   ;
  input                                           std__pe14__lane2_strm0_data_valid  ;

  output                                          pe14__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane2_strm1_data_mask   ;
  input                                           std__pe14__lane2_strm1_data_valid  ;

  output                                          pe14__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane3_strm0_data_mask   ;
  input                                           std__pe14__lane3_strm0_data_valid  ;

  output                                          pe14__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane3_strm1_data_mask   ;
  input                                           std__pe14__lane3_strm1_data_valid  ;

  output                                          pe14__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane4_strm0_data_mask   ;
  input                                           std__pe14__lane4_strm0_data_valid  ;

  output                                          pe14__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane4_strm1_data_mask   ;
  input                                           std__pe14__lane4_strm1_data_valid  ;

  output                                          pe14__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane5_strm0_data_mask   ;
  input                                           std__pe14__lane5_strm0_data_valid  ;

  output                                          pe14__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane5_strm1_data_mask   ;
  input                                           std__pe14__lane5_strm1_data_valid  ;

  output                                          pe14__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane6_strm0_data_mask   ;
  input                                           std__pe14__lane6_strm0_data_valid  ;

  output                                          pe14__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane6_strm1_data_mask   ;
  input                                           std__pe14__lane6_strm1_data_valid  ;

  output                                          pe14__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane7_strm0_data_mask   ;
  input                                           std__pe14__lane7_strm0_data_valid  ;

  output                                          pe14__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane7_strm1_data_mask   ;
  input                                           std__pe14__lane7_strm1_data_valid  ;

  output                                          pe14__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane8_strm0_data_mask   ;
  input                                           std__pe14__lane8_strm0_data_valid  ;

  output                                          pe14__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane8_strm1_data_mask   ;
  input                                           std__pe14__lane8_strm1_data_valid  ;

  output                                          pe14__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane9_strm0_data_mask   ;
  input                                           std__pe14__lane9_strm0_data_valid  ;

  output                                          pe14__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane9_strm1_data_mask   ;
  input                                           std__pe14__lane9_strm1_data_valid  ;

  output                                          pe14__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane10_strm0_data_mask   ;
  input                                           std__pe14__lane10_strm0_data_valid  ;

  output                                          pe14__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane10_strm1_data_mask   ;
  input                                           std__pe14__lane10_strm1_data_valid  ;

  output                                          pe14__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane11_strm0_data_mask   ;
  input                                           std__pe14__lane11_strm0_data_valid  ;

  output                                          pe14__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane11_strm1_data_mask   ;
  input                                           std__pe14__lane11_strm1_data_valid  ;

  output                                          pe14__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane12_strm0_data_mask   ;
  input                                           std__pe14__lane12_strm0_data_valid  ;

  output                                          pe14__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane12_strm1_data_mask   ;
  input                                           std__pe14__lane12_strm1_data_valid  ;

  output                                          pe14__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane13_strm0_data_mask   ;
  input                                           std__pe14__lane13_strm0_data_valid  ;

  output                                          pe14__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane13_strm1_data_mask   ;
  input                                           std__pe14__lane13_strm1_data_valid  ;

  output                                          pe14__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane14_strm0_data_mask   ;
  input                                           std__pe14__lane14_strm0_data_valid  ;

  output                                          pe14__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane14_strm1_data_mask   ;
  input                                           std__pe14__lane14_strm1_data_valid  ;

  output                                          pe14__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane15_strm0_data_mask   ;
  input                                           std__pe14__lane15_strm0_data_valid  ;

  output                                          pe14__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane15_strm1_data_mask   ;
  input                                           std__pe14__lane15_strm1_data_valid  ;

  output                                          pe14__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane16_strm0_data_mask   ;
  input                                           std__pe14__lane16_strm0_data_valid  ;

  output                                          pe14__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane16_strm1_data_mask   ;
  input                                           std__pe14__lane16_strm1_data_valid  ;

  output                                          pe14__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane17_strm0_data_mask   ;
  input                                           std__pe14__lane17_strm0_data_valid  ;

  output                                          pe14__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane17_strm1_data_mask   ;
  input                                           std__pe14__lane17_strm1_data_valid  ;

  output                                          pe14__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane18_strm0_data_mask   ;
  input                                           std__pe14__lane18_strm0_data_valid  ;

  output                                          pe14__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane18_strm1_data_mask   ;
  input                                           std__pe14__lane18_strm1_data_valid  ;

  output                                          pe14__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane19_strm0_data_mask   ;
  input                                           std__pe14__lane19_strm0_data_valid  ;

  output                                          pe14__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane19_strm1_data_mask   ;
  input                                           std__pe14__lane19_strm1_data_valid  ;

  output                                          pe14__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane20_strm0_data_mask   ;
  input                                           std__pe14__lane20_strm0_data_valid  ;

  output                                          pe14__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane20_strm1_data_mask   ;
  input                                           std__pe14__lane20_strm1_data_valid  ;

  output                                          pe14__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane21_strm0_data_mask   ;
  input                                           std__pe14__lane21_strm0_data_valid  ;

  output                                          pe14__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane21_strm1_data_mask   ;
  input                                           std__pe14__lane21_strm1_data_valid  ;

  output                                          pe14__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane22_strm0_data_mask   ;
  input                                           std__pe14__lane22_strm0_data_valid  ;

  output                                          pe14__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane22_strm1_data_mask   ;
  input                                           std__pe14__lane22_strm1_data_valid  ;

  output                                          pe14__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane23_strm0_data_mask   ;
  input                                           std__pe14__lane23_strm0_data_valid  ;

  output                                          pe14__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane23_strm1_data_mask   ;
  input                                           std__pe14__lane23_strm1_data_valid  ;

  output                                          pe14__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane24_strm0_data_mask   ;
  input                                           std__pe14__lane24_strm0_data_valid  ;

  output                                          pe14__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane24_strm1_data_mask   ;
  input                                           std__pe14__lane24_strm1_data_valid  ;

  output                                          pe14__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane25_strm0_data_mask   ;
  input                                           std__pe14__lane25_strm0_data_valid  ;

  output                                          pe14__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane25_strm1_data_mask   ;
  input                                           std__pe14__lane25_strm1_data_valid  ;

  output                                          pe14__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane26_strm0_data_mask   ;
  input                                           std__pe14__lane26_strm0_data_valid  ;

  output                                          pe14__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane26_strm1_data_mask   ;
  input                                           std__pe14__lane26_strm1_data_valid  ;

  output                                          pe14__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane27_strm0_data_mask   ;
  input                                           std__pe14__lane27_strm0_data_valid  ;

  output                                          pe14__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane27_strm1_data_mask   ;
  input                                           std__pe14__lane27_strm1_data_valid  ;

  output                                          pe14__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane28_strm0_data_mask   ;
  input                                           std__pe14__lane28_strm0_data_valid  ;

  output                                          pe14__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane28_strm1_data_mask   ;
  input                                           std__pe14__lane28_strm1_data_valid  ;

  output                                          pe14__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane29_strm0_data_mask   ;
  input                                           std__pe14__lane29_strm0_data_valid  ;

  output                                          pe14__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane29_strm1_data_mask   ;
  input                                           std__pe14__lane29_strm1_data_valid  ;

  output                                          pe14__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane30_strm0_data_mask   ;
  input                                           std__pe14__lane30_strm0_data_valid  ;

  output                                          pe14__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane30_strm1_data_mask   ;
  input                                           std__pe14__lane30_strm1_data_valid  ;

  output                                          pe14__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane31_strm0_data_mask   ;
  input                                           std__pe14__lane31_strm0_data_valid  ;

  output                                          pe14__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe14__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe14__lane31_strm1_data_mask   ;
  input                                           std__pe14__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe15__peId                ;
  input                                         sys__pe15__allSynchronized     ;
  output                                        pe15__sys__thisSynchronized    ;
  output                                        pe15__sys__ready               ;
  output                                        pe15__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe15__oob_cntl            ;
  input                                         std__pe15__oob_valid           ;
  output                                        pe15__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe15__oob_type            ;
  output                                          pe15__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane0_strm0_data_mask   ;
  input                                           std__pe15__lane0_strm0_data_valid  ;

  output                                          pe15__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane0_strm1_data_mask   ;
  input                                           std__pe15__lane0_strm1_data_valid  ;

  output                                          pe15__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane1_strm0_data_mask   ;
  input                                           std__pe15__lane1_strm0_data_valid  ;

  output                                          pe15__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane1_strm1_data_mask   ;
  input                                           std__pe15__lane1_strm1_data_valid  ;

  output                                          pe15__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane2_strm0_data_mask   ;
  input                                           std__pe15__lane2_strm0_data_valid  ;

  output                                          pe15__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane2_strm1_data_mask   ;
  input                                           std__pe15__lane2_strm1_data_valid  ;

  output                                          pe15__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane3_strm0_data_mask   ;
  input                                           std__pe15__lane3_strm0_data_valid  ;

  output                                          pe15__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane3_strm1_data_mask   ;
  input                                           std__pe15__lane3_strm1_data_valid  ;

  output                                          pe15__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane4_strm0_data_mask   ;
  input                                           std__pe15__lane4_strm0_data_valid  ;

  output                                          pe15__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane4_strm1_data_mask   ;
  input                                           std__pe15__lane4_strm1_data_valid  ;

  output                                          pe15__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane5_strm0_data_mask   ;
  input                                           std__pe15__lane5_strm0_data_valid  ;

  output                                          pe15__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane5_strm1_data_mask   ;
  input                                           std__pe15__lane5_strm1_data_valid  ;

  output                                          pe15__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane6_strm0_data_mask   ;
  input                                           std__pe15__lane6_strm0_data_valid  ;

  output                                          pe15__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane6_strm1_data_mask   ;
  input                                           std__pe15__lane6_strm1_data_valid  ;

  output                                          pe15__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane7_strm0_data_mask   ;
  input                                           std__pe15__lane7_strm0_data_valid  ;

  output                                          pe15__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane7_strm1_data_mask   ;
  input                                           std__pe15__lane7_strm1_data_valid  ;

  output                                          pe15__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane8_strm0_data_mask   ;
  input                                           std__pe15__lane8_strm0_data_valid  ;

  output                                          pe15__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane8_strm1_data_mask   ;
  input                                           std__pe15__lane8_strm1_data_valid  ;

  output                                          pe15__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane9_strm0_data_mask   ;
  input                                           std__pe15__lane9_strm0_data_valid  ;

  output                                          pe15__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane9_strm1_data_mask   ;
  input                                           std__pe15__lane9_strm1_data_valid  ;

  output                                          pe15__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane10_strm0_data_mask   ;
  input                                           std__pe15__lane10_strm0_data_valid  ;

  output                                          pe15__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane10_strm1_data_mask   ;
  input                                           std__pe15__lane10_strm1_data_valid  ;

  output                                          pe15__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane11_strm0_data_mask   ;
  input                                           std__pe15__lane11_strm0_data_valid  ;

  output                                          pe15__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane11_strm1_data_mask   ;
  input                                           std__pe15__lane11_strm1_data_valid  ;

  output                                          pe15__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane12_strm0_data_mask   ;
  input                                           std__pe15__lane12_strm0_data_valid  ;

  output                                          pe15__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane12_strm1_data_mask   ;
  input                                           std__pe15__lane12_strm1_data_valid  ;

  output                                          pe15__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane13_strm0_data_mask   ;
  input                                           std__pe15__lane13_strm0_data_valid  ;

  output                                          pe15__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane13_strm1_data_mask   ;
  input                                           std__pe15__lane13_strm1_data_valid  ;

  output                                          pe15__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane14_strm0_data_mask   ;
  input                                           std__pe15__lane14_strm0_data_valid  ;

  output                                          pe15__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane14_strm1_data_mask   ;
  input                                           std__pe15__lane14_strm1_data_valid  ;

  output                                          pe15__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane15_strm0_data_mask   ;
  input                                           std__pe15__lane15_strm0_data_valid  ;

  output                                          pe15__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane15_strm1_data_mask   ;
  input                                           std__pe15__lane15_strm1_data_valid  ;

  output                                          pe15__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane16_strm0_data_mask   ;
  input                                           std__pe15__lane16_strm0_data_valid  ;

  output                                          pe15__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane16_strm1_data_mask   ;
  input                                           std__pe15__lane16_strm1_data_valid  ;

  output                                          pe15__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane17_strm0_data_mask   ;
  input                                           std__pe15__lane17_strm0_data_valid  ;

  output                                          pe15__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane17_strm1_data_mask   ;
  input                                           std__pe15__lane17_strm1_data_valid  ;

  output                                          pe15__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane18_strm0_data_mask   ;
  input                                           std__pe15__lane18_strm0_data_valid  ;

  output                                          pe15__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane18_strm1_data_mask   ;
  input                                           std__pe15__lane18_strm1_data_valid  ;

  output                                          pe15__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane19_strm0_data_mask   ;
  input                                           std__pe15__lane19_strm0_data_valid  ;

  output                                          pe15__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane19_strm1_data_mask   ;
  input                                           std__pe15__lane19_strm1_data_valid  ;

  output                                          pe15__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane20_strm0_data_mask   ;
  input                                           std__pe15__lane20_strm0_data_valid  ;

  output                                          pe15__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane20_strm1_data_mask   ;
  input                                           std__pe15__lane20_strm1_data_valid  ;

  output                                          pe15__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane21_strm0_data_mask   ;
  input                                           std__pe15__lane21_strm0_data_valid  ;

  output                                          pe15__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane21_strm1_data_mask   ;
  input                                           std__pe15__lane21_strm1_data_valid  ;

  output                                          pe15__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane22_strm0_data_mask   ;
  input                                           std__pe15__lane22_strm0_data_valid  ;

  output                                          pe15__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane22_strm1_data_mask   ;
  input                                           std__pe15__lane22_strm1_data_valid  ;

  output                                          pe15__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane23_strm0_data_mask   ;
  input                                           std__pe15__lane23_strm0_data_valid  ;

  output                                          pe15__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane23_strm1_data_mask   ;
  input                                           std__pe15__lane23_strm1_data_valid  ;

  output                                          pe15__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane24_strm0_data_mask   ;
  input                                           std__pe15__lane24_strm0_data_valid  ;

  output                                          pe15__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane24_strm1_data_mask   ;
  input                                           std__pe15__lane24_strm1_data_valid  ;

  output                                          pe15__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane25_strm0_data_mask   ;
  input                                           std__pe15__lane25_strm0_data_valid  ;

  output                                          pe15__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane25_strm1_data_mask   ;
  input                                           std__pe15__lane25_strm1_data_valid  ;

  output                                          pe15__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane26_strm0_data_mask   ;
  input                                           std__pe15__lane26_strm0_data_valid  ;

  output                                          pe15__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane26_strm1_data_mask   ;
  input                                           std__pe15__lane26_strm1_data_valid  ;

  output                                          pe15__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane27_strm0_data_mask   ;
  input                                           std__pe15__lane27_strm0_data_valid  ;

  output                                          pe15__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane27_strm1_data_mask   ;
  input                                           std__pe15__lane27_strm1_data_valid  ;

  output                                          pe15__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane28_strm0_data_mask   ;
  input                                           std__pe15__lane28_strm0_data_valid  ;

  output                                          pe15__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane28_strm1_data_mask   ;
  input                                           std__pe15__lane28_strm1_data_valid  ;

  output                                          pe15__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane29_strm0_data_mask   ;
  input                                           std__pe15__lane29_strm0_data_valid  ;

  output                                          pe15__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane29_strm1_data_mask   ;
  input                                           std__pe15__lane29_strm1_data_valid  ;

  output                                          pe15__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane30_strm0_data_mask   ;
  input                                           std__pe15__lane30_strm0_data_valid  ;

  output                                          pe15__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane30_strm1_data_mask   ;
  input                                           std__pe15__lane30_strm1_data_valid  ;

  output                                          pe15__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane31_strm0_data_mask   ;
  input                                           std__pe15__lane31_strm0_data_valid  ;

  output                                          pe15__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe15__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe15__lane31_strm1_data_mask   ;
  input                                           std__pe15__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe16__peId                ;
  input                                         sys__pe16__allSynchronized     ;
  output                                        pe16__sys__thisSynchronized    ;
  output                                        pe16__sys__ready               ;
  output                                        pe16__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe16__oob_cntl            ;
  input                                         std__pe16__oob_valid           ;
  output                                        pe16__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe16__oob_type            ;
  output                                          pe16__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane0_strm0_data_mask   ;
  input                                           std__pe16__lane0_strm0_data_valid  ;

  output                                          pe16__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane0_strm1_data_mask   ;
  input                                           std__pe16__lane0_strm1_data_valid  ;

  output                                          pe16__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane1_strm0_data_mask   ;
  input                                           std__pe16__lane1_strm0_data_valid  ;

  output                                          pe16__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane1_strm1_data_mask   ;
  input                                           std__pe16__lane1_strm1_data_valid  ;

  output                                          pe16__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane2_strm0_data_mask   ;
  input                                           std__pe16__lane2_strm0_data_valid  ;

  output                                          pe16__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane2_strm1_data_mask   ;
  input                                           std__pe16__lane2_strm1_data_valid  ;

  output                                          pe16__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane3_strm0_data_mask   ;
  input                                           std__pe16__lane3_strm0_data_valid  ;

  output                                          pe16__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane3_strm1_data_mask   ;
  input                                           std__pe16__lane3_strm1_data_valid  ;

  output                                          pe16__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane4_strm0_data_mask   ;
  input                                           std__pe16__lane4_strm0_data_valid  ;

  output                                          pe16__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane4_strm1_data_mask   ;
  input                                           std__pe16__lane4_strm1_data_valid  ;

  output                                          pe16__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane5_strm0_data_mask   ;
  input                                           std__pe16__lane5_strm0_data_valid  ;

  output                                          pe16__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane5_strm1_data_mask   ;
  input                                           std__pe16__lane5_strm1_data_valid  ;

  output                                          pe16__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane6_strm0_data_mask   ;
  input                                           std__pe16__lane6_strm0_data_valid  ;

  output                                          pe16__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane6_strm1_data_mask   ;
  input                                           std__pe16__lane6_strm1_data_valid  ;

  output                                          pe16__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane7_strm0_data_mask   ;
  input                                           std__pe16__lane7_strm0_data_valid  ;

  output                                          pe16__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane7_strm1_data_mask   ;
  input                                           std__pe16__lane7_strm1_data_valid  ;

  output                                          pe16__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane8_strm0_data_mask   ;
  input                                           std__pe16__lane8_strm0_data_valid  ;

  output                                          pe16__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane8_strm1_data_mask   ;
  input                                           std__pe16__lane8_strm1_data_valid  ;

  output                                          pe16__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane9_strm0_data_mask   ;
  input                                           std__pe16__lane9_strm0_data_valid  ;

  output                                          pe16__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane9_strm1_data_mask   ;
  input                                           std__pe16__lane9_strm1_data_valid  ;

  output                                          pe16__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane10_strm0_data_mask   ;
  input                                           std__pe16__lane10_strm0_data_valid  ;

  output                                          pe16__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane10_strm1_data_mask   ;
  input                                           std__pe16__lane10_strm1_data_valid  ;

  output                                          pe16__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane11_strm0_data_mask   ;
  input                                           std__pe16__lane11_strm0_data_valid  ;

  output                                          pe16__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane11_strm1_data_mask   ;
  input                                           std__pe16__lane11_strm1_data_valid  ;

  output                                          pe16__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane12_strm0_data_mask   ;
  input                                           std__pe16__lane12_strm0_data_valid  ;

  output                                          pe16__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane12_strm1_data_mask   ;
  input                                           std__pe16__lane12_strm1_data_valid  ;

  output                                          pe16__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane13_strm0_data_mask   ;
  input                                           std__pe16__lane13_strm0_data_valid  ;

  output                                          pe16__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane13_strm1_data_mask   ;
  input                                           std__pe16__lane13_strm1_data_valid  ;

  output                                          pe16__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane14_strm0_data_mask   ;
  input                                           std__pe16__lane14_strm0_data_valid  ;

  output                                          pe16__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane14_strm1_data_mask   ;
  input                                           std__pe16__lane14_strm1_data_valid  ;

  output                                          pe16__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane15_strm0_data_mask   ;
  input                                           std__pe16__lane15_strm0_data_valid  ;

  output                                          pe16__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane15_strm1_data_mask   ;
  input                                           std__pe16__lane15_strm1_data_valid  ;

  output                                          pe16__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane16_strm0_data_mask   ;
  input                                           std__pe16__lane16_strm0_data_valid  ;

  output                                          pe16__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane16_strm1_data_mask   ;
  input                                           std__pe16__lane16_strm1_data_valid  ;

  output                                          pe16__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane17_strm0_data_mask   ;
  input                                           std__pe16__lane17_strm0_data_valid  ;

  output                                          pe16__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane17_strm1_data_mask   ;
  input                                           std__pe16__lane17_strm1_data_valid  ;

  output                                          pe16__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane18_strm0_data_mask   ;
  input                                           std__pe16__lane18_strm0_data_valid  ;

  output                                          pe16__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane18_strm1_data_mask   ;
  input                                           std__pe16__lane18_strm1_data_valid  ;

  output                                          pe16__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane19_strm0_data_mask   ;
  input                                           std__pe16__lane19_strm0_data_valid  ;

  output                                          pe16__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane19_strm1_data_mask   ;
  input                                           std__pe16__lane19_strm1_data_valid  ;

  output                                          pe16__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane20_strm0_data_mask   ;
  input                                           std__pe16__lane20_strm0_data_valid  ;

  output                                          pe16__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane20_strm1_data_mask   ;
  input                                           std__pe16__lane20_strm1_data_valid  ;

  output                                          pe16__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane21_strm0_data_mask   ;
  input                                           std__pe16__lane21_strm0_data_valid  ;

  output                                          pe16__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane21_strm1_data_mask   ;
  input                                           std__pe16__lane21_strm1_data_valid  ;

  output                                          pe16__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane22_strm0_data_mask   ;
  input                                           std__pe16__lane22_strm0_data_valid  ;

  output                                          pe16__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane22_strm1_data_mask   ;
  input                                           std__pe16__lane22_strm1_data_valid  ;

  output                                          pe16__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane23_strm0_data_mask   ;
  input                                           std__pe16__lane23_strm0_data_valid  ;

  output                                          pe16__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane23_strm1_data_mask   ;
  input                                           std__pe16__lane23_strm1_data_valid  ;

  output                                          pe16__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane24_strm0_data_mask   ;
  input                                           std__pe16__lane24_strm0_data_valid  ;

  output                                          pe16__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane24_strm1_data_mask   ;
  input                                           std__pe16__lane24_strm1_data_valid  ;

  output                                          pe16__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane25_strm0_data_mask   ;
  input                                           std__pe16__lane25_strm0_data_valid  ;

  output                                          pe16__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane25_strm1_data_mask   ;
  input                                           std__pe16__lane25_strm1_data_valid  ;

  output                                          pe16__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane26_strm0_data_mask   ;
  input                                           std__pe16__lane26_strm0_data_valid  ;

  output                                          pe16__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane26_strm1_data_mask   ;
  input                                           std__pe16__lane26_strm1_data_valid  ;

  output                                          pe16__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane27_strm0_data_mask   ;
  input                                           std__pe16__lane27_strm0_data_valid  ;

  output                                          pe16__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane27_strm1_data_mask   ;
  input                                           std__pe16__lane27_strm1_data_valid  ;

  output                                          pe16__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane28_strm0_data_mask   ;
  input                                           std__pe16__lane28_strm0_data_valid  ;

  output                                          pe16__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane28_strm1_data_mask   ;
  input                                           std__pe16__lane28_strm1_data_valid  ;

  output                                          pe16__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane29_strm0_data_mask   ;
  input                                           std__pe16__lane29_strm0_data_valid  ;

  output                                          pe16__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane29_strm1_data_mask   ;
  input                                           std__pe16__lane29_strm1_data_valid  ;

  output                                          pe16__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane30_strm0_data_mask   ;
  input                                           std__pe16__lane30_strm0_data_valid  ;

  output                                          pe16__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane30_strm1_data_mask   ;
  input                                           std__pe16__lane30_strm1_data_valid  ;

  output                                          pe16__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane31_strm0_data_mask   ;
  input                                           std__pe16__lane31_strm0_data_valid  ;

  output                                          pe16__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe16__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe16__lane31_strm1_data_mask   ;
  input                                           std__pe16__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe17__peId                ;
  input                                         sys__pe17__allSynchronized     ;
  output                                        pe17__sys__thisSynchronized    ;
  output                                        pe17__sys__ready               ;
  output                                        pe17__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe17__oob_cntl            ;
  input                                         std__pe17__oob_valid           ;
  output                                        pe17__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe17__oob_type            ;
  output                                          pe17__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane0_strm0_data_mask   ;
  input                                           std__pe17__lane0_strm0_data_valid  ;

  output                                          pe17__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane0_strm1_data_mask   ;
  input                                           std__pe17__lane0_strm1_data_valid  ;

  output                                          pe17__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane1_strm0_data_mask   ;
  input                                           std__pe17__lane1_strm0_data_valid  ;

  output                                          pe17__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane1_strm1_data_mask   ;
  input                                           std__pe17__lane1_strm1_data_valid  ;

  output                                          pe17__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane2_strm0_data_mask   ;
  input                                           std__pe17__lane2_strm0_data_valid  ;

  output                                          pe17__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane2_strm1_data_mask   ;
  input                                           std__pe17__lane2_strm1_data_valid  ;

  output                                          pe17__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane3_strm0_data_mask   ;
  input                                           std__pe17__lane3_strm0_data_valid  ;

  output                                          pe17__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane3_strm1_data_mask   ;
  input                                           std__pe17__lane3_strm1_data_valid  ;

  output                                          pe17__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane4_strm0_data_mask   ;
  input                                           std__pe17__lane4_strm0_data_valid  ;

  output                                          pe17__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane4_strm1_data_mask   ;
  input                                           std__pe17__lane4_strm1_data_valid  ;

  output                                          pe17__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane5_strm0_data_mask   ;
  input                                           std__pe17__lane5_strm0_data_valid  ;

  output                                          pe17__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane5_strm1_data_mask   ;
  input                                           std__pe17__lane5_strm1_data_valid  ;

  output                                          pe17__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane6_strm0_data_mask   ;
  input                                           std__pe17__lane6_strm0_data_valid  ;

  output                                          pe17__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane6_strm1_data_mask   ;
  input                                           std__pe17__lane6_strm1_data_valid  ;

  output                                          pe17__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane7_strm0_data_mask   ;
  input                                           std__pe17__lane7_strm0_data_valid  ;

  output                                          pe17__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane7_strm1_data_mask   ;
  input                                           std__pe17__lane7_strm1_data_valid  ;

  output                                          pe17__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane8_strm0_data_mask   ;
  input                                           std__pe17__lane8_strm0_data_valid  ;

  output                                          pe17__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane8_strm1_data_mask   ;
  input                                           std__pe17__lane8_strm1_data_valid  ;

  output                                          pe17__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane9_strm0_data_mask   ;
  input                                           std__pe17__lane9_strm0_data_valid  ;

  output                                          pe17__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane9_strm1_data_mask   ;
  input                                           std__pe17__lane9_strm1_data_valid  ;

  output                                          pe17__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane10_strm0_data_mask   ;
  input                                           std__pe17__lane10_strm0_data_valid  ;

  output                                          pe17__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane10_strm1_data_mask   ;
  input                                           std__pe17__lane10_strm1_data_valid  ;

  output                                          pe17__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane11_strm0_data_mask   ;
  input                                           std__pe17__lane11_strm0_data_valid  ;

  output                                          pe17__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane11_strm1_data_mask   ;
  input                                           std__pe17__lane11_strm1_data_valid  ;

  output                                          pe17__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane12_strm0_data_mask   ;
  input                                           std__pe17__lane12_strm0_data_valid  ;

  output                                          pe17__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane12_strm1_data_mask   ;
  input                                           std__pe17__lane12_strm1_data_valid  ;

  output                                          pe17__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane13_strm0_data_mask   ;
  input                                           std__pe17__lane13_strm0_data_valid  ;

  output                                          pe17__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane13_strm1_data_mask   ;
  input                                           std__pe17__lane13_strm1_data_valid  ;

  output                                          pe17__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane14_strm0_data_mask   ;
  input                                           std__pe17__lane14_strm0_data_valid  ;

  output                                          pe17__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane14_strm1_data_mask   ;
  input                                           std__pe17__lane14_strm1_data_valid  ;

  output                                          pe17__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane15_strm0_data_mask   ;
  input                                           std__pe17__lane15_strm0_data_valid  ;

  output                                          pe17__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane15_strm1_data_mask   ;
  input                                           std__pe17__lane15_strm1_data_valid  ;

  output                                          pe17__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane16_strm0_data_mask   ;
  input                                           std__pe17__lane16_strm0_data_valid  ;

  output                                          pe17__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane16_strm1_data_mask   ;
  input                                           std__pe17__lane16_strm1_data_valid  ;

  output                                          pe17__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane17_strm0_data_mask   ;
  input                                           std__pe17__lane17_strm0_data_valid  ;

  output                                          pe17__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane17_strm1_data_mask   ;
  input                                           std__pe17__lane17_strm1_data_valid  ;

  output                                          pe17__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane18_strm0_data_mask   ;
  input                                           std__pe17__lane18_strm0_data_valid  ;

  output                                          pe17__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane18_strm1_data_mask   ;
  input                                           std__pe17__lane18_strm1_data_valid  ;

  output                                          pe17__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane19_strm0_data_mask   ;
  input                                           std__pe17__lane19_strm0_data_valid  ;

  output                                          pe17__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane19_strm1_data_mask   ;
  input                                           std__pe17__lane19_strm1_data_valid  ;

  output                                          pe17__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane20_strm0_data_mask   ;
  input                                           std__pe17__lane20_strm0_data_valid  ;

  output                                          pe17__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane20_strm1_data_mask   ;
  input                                           std__pe17__lane20_strm1_data_valid  ;

  output                                          pe17__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane21_strm0_data_mask   ;
  input                                           std__pe17__lane21_strm0_data_valid  ;

  output                                          pe17__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane21_strm1_data_mask   ;
  input                                           std__pe17__lane21_strm1_data_valid  ;

  output                                          pe17__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane22_strm0_data_mask   ;
  input                                           std__pe17__lane22_strm0_data_valid  ;

  output                                          pe17__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane22_strm1_data_mask   ;
  input                                           std__pe17__lane22_strm1_data_valid  ;

  output                                          pe17__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane23_strm0_data_mask   ;
  input                                           std__pe17__lane23_strm0_data_valid  ;

  output                                          pe17__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane23_strm1_data_mask   ;
  input                                           std__pe17__lane23_strm1_data_valid  ;

  output                                          pe17__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane24_strm0_data_mask   ;
  input                                           std__pe17__lane24_strm0_data_valid  ;

  output                                          pe17__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane24_strm1_data_mask   ;
  input                                           std__pe17__lane24_strm1_data_valid  ;

  output                                          pe17__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane25_strm0_data_mask   ;
  input                                           std__pe17__lane25_strm0_data_valid  ;

  output                                          pe17__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane25_strm1_data_mask   ;
  input                                           std__pe17__lane25_strm1_data_valid  ;

  output                                          pe17__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane26_strm0_data_mask   ;
  input                                           std__pe17__lane26_strm0_data_valid  ;

  output                                          pe17__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane26_strm1_data_mask   ;
  input                                           std__pe17__lane26_strm1_data_valid  ;

  output                                          pe17__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane27_strm0_data_mask   ;
  input                                           std__pe17__lane27_strm0_data_valid  ;

  output                                          pe17__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane27_strm1_data_mask   ;
  input                                           std__pe17__lane27_strm1_data_valid  ;

  output                                          pe17__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane28_strm0_data_mask   ;
  input                                           std__pe17__lane28_strm0_data_valid  ;

  output                                          pe17__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane28_strm1_data_mask   ;
  input                                           std__pe17__lane28_strm1_data_valid  ;

  output                                          pe17__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane29_strm0_data_mask   ;
  input                                           std__pe17__lane29_strm0_data_valid  ;

  output                                          pe17__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane29_strm1_data_mask   ;
  input                                           std__pe17__lane29_strm1_data_valid  ;

  output                                          pe17__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane30_strm0_data_mask   ;
  input                                           std__pe17__lane30_strm0_data_valid  ;

  output                                          pe17__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane30_strm1_data_mask   ;
  input                                           std__pe17__lane30_strm1_data_valid  ;

  output                                          pe17__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane31_strm0_data_mask   ;
  input                                           std__pe17__lane31_strm0_data_valid  ;

  output                                          pe17__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe17__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe17__lane31_strm1_data_mask   ;
  input                                           std__pe17__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe18__peId                ;
  input                                         sys__pe18__allSynchronized     ;
  output                                        pe18__sys__thisSynchronized    ;
  output                                        pe18__sys__ready               ;
  output                                        pe18__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe18__oob_cntl            ;
  input                                         std__pe18__oob_valid           ;
  output                                        pe18__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe18__oob_type            ;
  output                                          pe18__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane0_strm0_data_mask   ;
  input                                           std__pe18__lane0_strm0_data_valid  ;

  output                                          pe18__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane0_strm1_data_mask   ;
  input                                           std__pe18__lane0_strm1_data_valid  ;

  output                                          pe18__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane1_strm0_data_mask   ;
  input                                           std__pe18__lane1_strm0_data_valid  ;

  output                                          pe18__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane1_strm1_data_mask   ;
  input                                           std__pe18__lane1_strm1_data_valid  ;

  output                                          pe18__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane2_strm0_data_mask   ;
  input                                           std__pe18__lane2_strm0_data_valid  ;

  output                                          pe18__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane2_strm1_data_mask   ;
  input                                           std__pe18__lane2_strm1_data_valid  ;

  output                                          pe18__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane3_strm0_data_mask   ;
  input                                           std__pe18__lane3_strm0_data_valid  ;

  output                                          pe18__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane3_strm1_data_mask   ;
  input                                           std__pe18__lane3_strm1_data_valid  ;

  output                                          pe18__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane4_strm0_data_mask   ;
  input                                           std__pe18__lane4_strm0_data_valid  ;

  output                                          pe18__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane4_strm1_data_mask   ;
  input                                           std__pe18__lane4_strm1_data_valid  ;

  output                                          pe18__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane5_strm0_data_mask   ;
  input                                           std__pe18__lane5_strm0_data_valid  ;

  output                                          pe18__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane5_strm1_data_mask   ;
  input                                           std__pe18__lane5_strm1_data_valid  ;

  output                                          pe18__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane6_strm0_data_mask   ;
  input                                           std__pe18__lane6_strm0_data_valid  ;

  output                                          pe18__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane6_strm1_data_mask   ;
  input                                           std__pe18__lane6_strm1_data_valid  ;

  output                                          pe18__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane7_strm0_data_mask   ;
  input                                           std__pe18__lane7_strm0_data_valid  ;

  output                                          pe18__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane7_strm1_data_mask   ;
  input                                           std__pe18__lane7_strm1_data_valid  ;

  output                                          pe18__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane8_strm0_data_mask   ;
  input                                           std__pe18__lane8_strm0_data_valid  ;

  output                                          pe18__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane8_strm1_data_mask   ;
  input                                           std__pe18__lane8_strm1_data_valid  ;

  output                                          pe18__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane9_strm0_data_mask   ;
  input                                           std__pe18__lane9_strm0_data_valid  ;

  output                                          pe18__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane9_strm1_data_mask   ;
  input                                           std__pe18__lane9_strm1_data_valid  ;

  output                                          pe18__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane10_strm0_data_mask   ;
  input                                           std__pe18__lane10_strm0_data_valid  ;

  output                                          pe18__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane10_strm1_data_mask   ;
  input                                           std__pe18__lane10_strm1_data_valid  ;

  output                                          pe18__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane11_strm0_data_mask   ;
  input                                           std__pe18__lane11_strm0_data_valid  ;

  output                                          pe18__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane11_strm1_data_mask   ;
  input                                           std__pe18__lane11_strm1_data_valid  ;

  output                                          pe18__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane12_strm0_data_mask   ;
  input                                           std__pe18__lane12_strm0_data_valid  ;

  output                                          pe18__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane12_strm1_data_mask   ;
  input                                           std__pe18__lane12_strm1_data_valid  ;

  output                                          pe18__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane13_strm0_data_mask   ;
  input                                           std__pe18__lane13_strm0_data_valid  ;

  output                                          pe18__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane13_strm1_data_mask   ;
  input                                           std__pe18__lane13_strm1_data_valid  ;

  output                                          pe18__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane14_strm0_data_mask   ;
  input                                           std__pe18__lane14_strm0_data_valid  ;

  output                                          pe18__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane14_strm1_data_mask   ;
  input                                           std__pe18__lane14_strm1_data_valid  ;

  output                                          pe18__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane15_strm0_data_mask   ;
  input                                           std__pe18__lane15_strm0_data_valid  ;

  output                                          pe18__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane15_strm1_data_mask   ;
  input                                           std__pe18__lane15_strm1_data_valid  ;

  output                                          pe18__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane16_strm0_data_mask   ;
  input                                           std__pe18__lane16_strm0_data_valid  ;

  output                                          pe18__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane16_strm1_data_mask   ;
  input                                           std__pe18__lane16_strm1_data_valid  ;

  output                                          pe18__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane17_strm0_data_mask   ;
  input                                           std__pe18__lane17_strm0_data_valid  ;

  output                                          pe18__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane17_strm1_data_mask   ;
  input                                           std__pe18__lane17_strm1_data_valid  ;

  output                                          pe18__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane18_strm0_data_mask   ;
  input                                           std__pe18__lane18_strm0_data_valid  ;

  output                                          pe18__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane18_strm1_data_mask   ;
  input                                           std__pe18__lane18_strm1_data_valid  ;

  output                                          pe18__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane19_strm0_data_mask   ;
  input                                           std__pe18__lane19_strm0_data_valid  ;

  output                                          pe18__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane19_strm1_data_mask   ;
  input                                           std__pe18__lane19_strm1_data_valid  ;

  output                                          pe18__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane20_strm0_data_mask   ;
  input                                           std__pe18__lane20_strm0_data_valid  ;

  output                                          pe18__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane20_strm1_data_mask   ;
  input                                           std__pe18__lane20_strm1_data_valid  ;

  output                                          pe18__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane21_strm0_data_mask   ;
  input                                           std__pe18__lane21_strm0_data_valid  ;

  output                                          pe18__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane21_strm1_data_mask   ;
  input                                           std__pe18__lane21_strm1_data_valid  ;

  output                                          pe18__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane22_strm0_data_mask   ;
  input                                           std__pe18__lane22_strm0_data_valid  ;

  output                                          pe18__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane22_strm1_data_mask   ;
  input                                           std__pe18__lane22_strm1_data_valid  ;

  output                                          pe18__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane23_strm0_data_mask   ;
  input                                           std__pe18__lane23_strm0_data_valid  ;

  output                                          pe18__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane23_strm1_data_mask   ;
  input                                           std__pe18__lane23_strm1_data_valid  ;

  output                                          pe18__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane24_strm0_data_mask   ;
  input                                           std__pe18__lane24_strm0_data_valid  ;

  output                                          pe18__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane24_strm1_data_mask   ;
  input                                           std__pe18__lane24_strm1_data_valid  ;

  output                                          pe18__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane25_strm0_data_mask   ;
  input                                           std__pe18__lane25_strm0_data_valid  ;

  output                                          pe18__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane25_strm1_data_mask   ;
  input                                           std__pe18__lane25_strm1_data_valid  ;

  output                                          pe18__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane26_strm0_data_mask   ;
  input                                           std__pe18__lane26_strm0_data_valid  ;

  output                                          pe18__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane26_strm1_data_mask   ;
  input                                           std__pe18__lane26_strm1_data_valid  ;

  output                                          pe18__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane27_strm0_data_mask   ;
  input                                           std__pe18__lane27_strm0_data_valid  ;

  output                                          pe18__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane27_strm1_data_mask   ;
  input                                           std__pe18__lane27_strm1_data_valid  ;

  output                                          pe18__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane28_strm0_data_mask   ;
  input                                           std__pe18__lane28_strm0_data_valid  ;

  output                                          pe18__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane28_strm1_data_mask   ;
  input                                           std__pe18__lane28_strm1_data_valid  ;

  output                                          pe18__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane29_strm0_data_mask   ;
  input                                           std__pe18__lane29_strm0_data_valid  ;

  output                                          pe18__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane29_strm1_data_mask   ;
  input                                           std__pe18__lane29_strm1_data_valid  ;

  output                                          pe18__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane30_strm0_data_mask   ;
  input                                           std__pe18__lane30_strm0_data_valid  ;

  output                                          pe18__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane30_strm1_data_mask   ;
  input                                           std__pe18__lane30_strm1_data_valid  ;

  output                                          pe18__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane31_strm0_data_mask   ;
  input                                           std__pe18__lane31_strm0_data_valid  ;

  output                                          pe18__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe18__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe18__lane31_strm1_data_mask   ;
  input                                           std__pe18__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe19__peId                ;
  input                                         sys__pe19__allSynchronized     ;
  output                                        pe19__sys__thisSynchronized    ;
  output                                        pe19__sys__ready               ;
  output                                        pe19__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe19__oob_cntl            ;
  input                                         std__pe19__oob_valid           ;
  output                                        pe19__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe19__oob_type            ;
  output                                          pe19__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane0_strm0_data_mask   ;
  input                                           std__pe19__lane0_strm0_data_valid  ;

  output                                          pe19__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane0_strm1_data_mask   ;
  input                                           std__pe19__lane0_strm1_data_valid  ;

  output                                          pe19__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane1_strm0_data_mask   ;
  input                                           std__pe19__lane1_strm0_data_valid  ;

  output                                          pe19__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane1_strm1_data_mask   ;
  input                                           std__pe19__lane1_strm1_data_valid  ;

  output                                          pe19__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane2_strm0_data_mask   ;
  input                                           std__pe19__lane2_strm0_data_valid  ;

  output                                          pe19__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane2_strm1_data_mask   ;
  input                                           std__pe19__lane2_strm1_data_valid  ;

  output                                          pe19__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane3_strm0_data_mask   ;
  input                                           std__pe19__lane3_strm0_data_valid  ;

  output                                          pe19__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane3_strm1_data_mask   ;
  input                                           std__pe19__lane3_strm1_data_valid  ;

  output                                          pe19__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane4_strm0_data_mask   ;
  input                                           std__pe19__lane4_strm0_data_valid  ;

  output                                          pe19__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane4_strm1_data_mask   ;
  input                                           std__pe19__lane4_strm1_data_valid  ;

  output                                          pe19__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane5_strm0_data_mask   ;
  input                                           std__pe19__lane5_strm0_data_valid  ;

  output                                          pe19__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane5_strm1_data_mask   ;
  input                                           std__pe19__lane5_strm1_data_valid  ;

  output                                          pe19__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane6_strm0_data_mask   ;
  input                                           std__pe19__lane6_strm0_data_valid  ;

  output                                          pe19__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane6_strm1_data_mask   ;
  input                                           std__pe19__lane6_strm1_data_valid  ;

  output                                          pe19__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane7_strm0_data_mask   ;
  input                                           std__pe19__lane7_strm0_data_valid  ;

  output                                          pe19__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane7_strm1_data_mask   ;
  input                                           std__pe19__lane7_strm1_data_valid  ;

  output                                          pe19__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane8_strm0_data_mask   ;
  input                                           std__pe19__lane8_strm0_data_valid  ;

  output                                          pe19__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane8_strm1_data_mask   ;
  input                                           std__pe19__lane8_strm1_data_valid  ;

  output                                          pe19__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane9_strm0_data_mask   ;
  input                                           std__pe19__lane9_strm0_data_valid  ;

  output                                          pe19__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane9_strm1_data_mask   ;
  input                                           std__pe19__lane9_strm1_data_valid  ;

  output                                          pe19__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane10_strm0_data_mask   ;
  input                                           std__pe19__lane10_strm0_data_valid  ;

  output                                          pe19__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane10_strm1_data_mask   ;
  input                                           std__pe19__lane10_strm1_data_valid  ;

  output                                          pe19__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane11_strm0_data_mask   ;
  input                                           std__pe19__lane11_strm0_data_valid  ;

  output                                          pe19__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane11_strm1_data_mask   ;
  input                                           std__pe19__lane11_strm1_data_valid  ;

  output                                          pe19__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane12_strm0_data_mask   ;
  input                                           std__pe19__lane12_strm0_data_valid  ;

  output                                          pe19__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane12_strm1_data_mask   ;
  input                                           std__pe19__lane12_strm1_data_valid  ;

  output                                          pe19__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane13_strm0_data_mask   ;
  input                                           std__pe19__lane13_strm0_data_valid  ;

  output                                          pe19__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane13_strm1_data_mask   ;
  input                                           std__pe19__lane13_strm1_data_valid  ;

  output                                          pe19__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane14_strm0_data_mask   ;
  input                                           std__pe19__lane14_strm0_data_valid  ;

  output                                          pe19__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane14_strm1_data_mask   ;
  input                                           std__pe19__lane14_strm1_data_valid  ;

  output                                          pe19__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane15_strm0_data_mask   ;
  input                                           std__pe19__lane15_strm0_data_valid  ;

  output                                          pe19__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane15_strm1_data_mask   ;
  input                                           std__pe19__lane15_strm1_data_valid  ;

  output                                          pe19__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane16_strm0_data_mask   ;
  input                                           std__pe19__lane16_strm0_data_valid  ;

  output                                          pe19__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane16_strm1_data_mask   ;
  input                                           std__pe19__lane16_strm1_data_valid  ;

  output                                          pe19__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane17_strm0_data_mask   ;
  input                                           std__pe19__lane17_strm0_data_valid  ;

  output                                          pe19__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane17_strm1_data_mask   ;
  input                                           std__pe19__lane17_strm1_data_valid  ;

  output                                          pe19__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane18_strm0_data_mask   ;
  input                                           std__pe19__lane18_strm0_data_valid  ;

  output                                          pe19__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane18_strm1_data_mask   ;
  input                                           std__pe19__lane18_strm1_data_valid  ;

  output                                          pe19__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane19_strm0_data_mask   ;
  input                                           std__pe19__lane19_strm0_data_valid  ;

  output                                          pe19__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane19_strm1_data_mask   ;
  input                                           std__pe19__lane19_strm1_data_valid  ;

  output                                          pe19__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane20_strm0_data_mask   ;
  input                                           std__pe19__lane20_strm0_data_valid  ;

  output                                          pe19__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane20_strm1_data_mask   ;
  input                                           std__pe19__lane20_strm1_data_valid  ;

  output                                          pe19__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane21_strm0_data_mask   ;
  input                                           std__pe19__lane21_strm0_data_valid  ;

  output                                          pe19__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane21_strm1_data_mask   ;
  input                                           std__pe19__lane21_strm1_data_valid  ;

  output                                          pe19__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane22_strm0_data_mask   ;
  input                                           std__pe19__lane22_strm0_data_valid  ;

  output                                          pe19__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane22_strm1_data_mask   ;
  input                                           std__pe19__lane22_strm1_data_valid  ;

  output                                          pe19__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane23_strm0_data_mask   ;
  input                                           std__pe19__lane23_strm0_data_valid  ;

  output                                          pe19__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane23_strm1_data_mask   ;
  input                                           std__pe19__lane23_strm1_data_valid  ;

  output                                          pe19__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane24_strm0_data_mask   ;
  input                                           std__pe19__lane24_strm0_data_valid  ;

  output                                          pe19__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane24_strm1_data_mask   ;
  input                                           std__pe19__lane24_strm1_data_valid  ;

  output                                          pe19__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane25_strm0_data_mask   ;
  input                                           std__pe19__lane25_strm0_data_valid  ;

  output                                          pe19__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane25_strm1_data_mask   ;
  input                                           std__pe19__lane25_strm1_data_valid  ;

  output                                          pe19__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane26_strm0_data_mask   ;
  input                                           std__pe19__lane26_strm0_data_valid  ;

  output                                          pe19__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane26_strm1_data_mask   ;
  input                                           std__pe19__lane26_strm1_data_valid  ;

  output                                          pe19__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane27_strm0_data_mask   ;
  input                                           std__pe19__lane27_strm0_data_valid  ;

  output                                          pe19__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane27_strm1_data_mask   ;
  input                                           std__pe19__lane27_strm1_data_valid  ;

  output                                          pe19__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane28_strm0_data_mask   ;
  input                                           std__pe19__lane28_strm0_data_valid  ;

  output                                          pe19__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane28_strm1_data_mask   ;
  input                                           std__pe19__lane28_strm1_data_valid  ;

  output                                          pe19__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane29_strm0_data_mask   ;
  input                                           std__pe19__lane29_strm0_data_valid  ;

  output                                          pe19__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane29_strm1_data_mask   ;
  input                                           std__pe19__lane29_strm1_data_valid  ;

  output                                          pe19__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane30_strm0_data_mask   ;
  input                                           std__pe19__lane30_strm0_data_valid  ;

  output                                          pe19__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane30_strm1_data_mask   ;
  input                                           std__pe19__lane30_strm1_data_valid  ;

  output                                          pe19__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane31_strm0_data_mask   ;
  input                                           std__pe19__lane31_strm0_data_valid  ;

  output                                          pe19__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe19__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe19__lane31_strm1_data_mask   ;
  input                                           std__pe19__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe20__peId                ;
  input                                         sys__pe20__allSynchronized     ;
  output                                        pe20__sys__thisSynchronized    ;
  output                                        pe20__sys__ready               ;
  output                                        pe20__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe20__oob_cntl            ;
  input                                         std__pe20__oob_valid           ;
  output                                        pe20__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe20__oob_type            ;
  output                                          pe20__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane0_strm0_data_mask   ;
  input                                           std__pe20__lane0_strm0_data_valid  ;

  output                                          pe20__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane0_strm1_data_mask   ;
  input                                           std__pe20__lane0_strm1_data_valid  ;

  output                                          pe20__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane1_strm0_data_mask   ;
  input                                           std__pe20__lane1_strm0_data_valid  ;

  output                                          pe20__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane1_strm1_data_mask   ;
  input                                           std__pe20__lane1_strm1_data_valid  ;

  output                                          pe20__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane2_strm0_data_mask   ;
  input                                           std__pe20__lane2_strm0_data_valid  ;

  output                                          pe20__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane2_strm1_data_mask   ;
  input                                           std__pe20__lane2_strm1_data_valid  ;

  output                                          pe20__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane3_strm0_data_mask   ;
  input                                           std__pe20__lane3_strm0_data_valid  ;

  output                                          pe20__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane3_strm1_data_mask   ;
  input                                           std__pe20__lane3_strm1_data_valid  ;

  output                                          pe20__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane4_strm0_data_mask   ;
  input                                           std__pe20__lane4_strm0_data_valid  ;

  output                                          pe20__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane4_strm1_data_mask   ;
  input                                           std__pe20__lane4_strm1_data_valid  ;

  output                                          pe20__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane5_strm0_data_mask   ;
  input                                           std__pe20__lane5_strm0_data_valid  ;

  output                                          pe20__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane5_strm1_data_mask   ;
  input                                           std__pe20__lane5_strm1_data_valid  ;

  output                                          pe20__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane6_strm0_data_mask   ;
  input                                           std__pe20__lane6_strm0_data_valid  ;

  output                                          pe20__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane6_strm1_data_mask   ;
  input                                           std__pe20__lane6_strm1_data_valid  ;

  output                                          pe20__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane7_strm0_data_mask   ;
  input                                           std__pe20__lane7_strm0_data_valid  ;

  output                                          pe20__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane7_strm1_data_mask   ;
  input                                           std__pe20__lane7_strm1_data_valid  ;

  output                                          pe20__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane8_strm0_data_mask   ;
  input                                           std__pe20__lane8_strm0_data_valid  ;

  output                                          pe20__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane8_strm1_data_mask   ;
  input                                           std__pe20__lane8_strm1_data_valid  ;

  output                                          pe20__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane9_strm0_data_mask   ;
  input                                           std__pe20__lane9_strm0_data_valid  ;

  output                                          pe20__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane9_strm1_data_mask   ;
  input                                           std__pe20__lane9_strm1_data_valid  ;

  output                                          pe20__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane10_strm0_data_mask   ;
  input                                           std__pe20__lane10_strm0_data_valid  ;

  output                                          pe20__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane10_strm1_data_mask   ;
  input                                           std__pe20__lane10_strm1_data_valid  ;

  output                                          pe20__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane11_strm0_data_mask   ;
  input                                           std__pe20__lane11_strm0_data_valid  ;

  output                                          pe20__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane11_strm1_data_mask   ;
  input                                           std__pe20__lane11_strm1_data_valid  ;

  output                                          pe20__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane12_strm0_data_mask   ;
  input                                           std__pe20__lane12_strm0_data_valid  ;

  output                                          pe20__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane12_strm1_data_mask   ;
  input                                           std__pe20__lane12_strm1_data_valid  ;

  output                                          pe20__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane13_strm0_data_mask   ;
  input                                           std__pe20__lane13_strm0_data_valid  ;

  output                                          pe20__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane13_strm1_data_mask   ;
  input                                           std__pe20__lane13_strm1_data_valid  ;

  output                                          pe20__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane14_strm0_data_mask   ;
  input                                           std__pe20__lane14_strm0_data_valid  ;

  output                                          pe20__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane14_strm1_data_mask   ;
  input                                           std__pe20__lane14_strm1_data_valid  ;

  output                                          pe20__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane15_strm0_data_mask   ;
  input                                           std__pe20__lane15_strm0_data_valid  ;

  output                                          pe20__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane15_strm1_data_mask   ;
  input                                           std__pe20__lane15_strm1_data_valid  ;

  output                                          pe20__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane16_strm0_data_mask   ;
  input                                           std__pe20__lane16_strm0_data_valid  ;

  output                                          pe20__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane16_strm1_data_mask   ;
  input                                           std__pe20__lane16_strm1_data_valid  ;

  output                                          pe20__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane17_strm0_data_mask   ;
  input                                           std__pe20__lane17_strm0_data_valid  ;

  output                                          pe20__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane17_strm1_data_mask   ;
  input                                           std__pe20__lane17_strm1_data_valid  ;

  output                                          pe20__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane18_strm0_data_mask   ;
  input                                           std__pe20__lane18_strm0_data_valid  ;

  output                                          pe20__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane18_strm1_data_mask   ;
  input                                           std__pe20__lane18_strm1_data_valid  ;

  output                                          pe20__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane19_strm0_data_mask   ;
  input                                           std__pe20__lane19_strm0_data_valid  ;

  output                                          pe20__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane19_strm1_data_mask   ;
  input                                           std__pe20__lane19_strm1_data_valid  ;

  output                                          pe20__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane20_strm0_data_mask   ;
  input                                           std__pe20__lane20_strm0_data_valid  ;

  output                                          pe20__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane20_strm1_data_mask   ;
  input                                           std__pe20__lane20_strm1_data_valid  ;

  output                                          pe20__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane21_strm0_data_mask   ;
  input                                           std__pe20__lane21_strm0_data_valid  ;

  output                                          pe20__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane21_strm1_data_mask   ;
  input                                           std__pe20__lane21_strm1_data_valid  ;

  output                                          pe20__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane22_strm0_data_mask   ;
  input                                           std__pe20__lane22_strm0_data_valid  ;

  output                                          pe20__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane22_strm1_data_mask   ;
  input                                           std__pe20__lane22_strm1_data_valid  ;

  output                                          pe20__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane23_strm0_data_mask   ;
  input                                           std__pe20__lane23_strm0_data_valid  ;

  output                                          pe20__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane23_strm1_data_mask   ;
  input                                           std__pe20__lane23_strm1_data_valid  ;

  output                                          pe20__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane24_strm0_data_mask   ;
  input                                           std__pe20__lane24_strm0_data_valid  ;

  output                                          pe20__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane24_strm1_data_mask   ;
  input                                           std__pe20__lane24_strm1_data_valid  ;

  output                                          pe20__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane25_strm0_data_mask   ;
  input                                           std__pe20__lane25_strm0_data_valid  ;

  output                                          pe20__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane25_strm1_data_mask   ;
  input                                           std__pe20__lane25_strm1_data_valid  ;

  output                                          pe20__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane26_strm0_data_mask   ;
  input                                           std__pe20__lane26_strm0_data_valid  ;

  output                                          pe20__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane26_strm1_data_mask   ;
  input                                           std__pe20__lane26_strm1_data_valid  ;

  output                                          pe20__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane27_strm0_data_mask   ;
  input                                           std__pe20__lane27_strm0_data_valid  ;

  output                                          pe20__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane27_strm1_data_mask   ;
  input                                           std__pe20__lane27_strm1_data_valid  ;

  output                                          pe20__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane28_strm0_data_mask   ;
  input                                           std__pe20__lane28_strm0_data_valid  ;

  output                                          pe20__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane28_strm1_data_mask   ;
  input                                           std__pe20__lane28_strm1_data_valid  ;

  output                                          pe20__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane29_strm0_data_mask   ;
  input                                           std__pe20__lane29_strm0_data_valid  ;

  output                                          pe20__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane29_strm1_data_mask   ;
  input                                           std__pe20__lane29_strm1_data_valid  ;

  output                                          pe20__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane30_strm0_data_mask   ;
  input                                           std__pe20__lane30_strm0_data_valid  ;

  output                                          pe20__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane30_strm1_data_mask   ;
  input                                           std__pe20__lane30_strm1_data_valid  ;

  output                                          pe20__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane31_strm0_data_mask   ;
  input                                           std__pe20__lane31_strm0_data_valid  ;

  output                                          pe20__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe20__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe20__lane31_strm1_data_mask   ;
  input                                           std__pe20__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe21__peId                ;
  input                                         sys__pe21__allSynchronized     ;
  output                                        pe21__sys__thisSynchronized    ;
  output                                        pe21__sys__ready               ;
  output                                        pe21__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe21__oob_cntl            ;
  input                                         std__pe21__oob_valid           ;
  output                                        pe21__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe21__oob_type            ;
  output                                          pe21__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane0_strm0_data_mask   ;
  input                                           std__pe21__lane0_strm0_data_valid  ;

  output                                          pe21__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane0_strm1_data_mask   ;
  input                                           std__pe21__lane0_strm1_data_valid  ;

  output                                          pe21__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane1_strm0_data_mask   ;
  input                                           std__pe21__lane1_strm0_data_valid  ;

  output                                          pe21__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane1_strm1_data_mask   ;
  input                                           std__pe21__lane1_strm1_data_valid  ;

  output                                          pe21__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane2_strm0_data_mask   ;
  input                                           std__pe21__lane2_strm0_data_valid  ;

  output                                          pe21__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane2_strm1_data_mask   ;
  input                                           std__pe21__lane2_strm1_data_valid  ;

  output                                          pe21__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane3_strm0_data_mask   ;
  input                                           std__pe21__lane3_strm0_data_valid  ;

  output                                          pe21__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane3_strm1_data_mask   ;
  input                                           std__pe21__lane3_strm1_data_valid  ;

  output                                          pe21__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane4_strm0_data_mask   ;
  input                                           std__pe21__lane4_strm0_data_valid  ;

  output                                          pe21__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane4_strm1_data_mask   ;
  input                                           std__pe21__lane4_strm1_data_valid  ;

  output                                          pe21__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane5_strm0_data_mask   ;
  input                                           std__pe21__lane5_strm0_data_valid  ;

  output                                          pe21__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane5_strm1_data_mask   ;
  input                                           std__pe21__lane5_strm1_data_valid  ;

  output                                          pe21__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane6_strm0_data_mask   ;
  input                                           std__pe21__lane6_strm0_data_valid  ;

  output                                          pe21__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane6_strm1_data_mask   ;
  input                                           std__pe21__lane6_strm1_data_valid  ;

  output                                          pe21__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane7_strm0_data_mask   ;
  input                                           std__pe21__lane7_strm0_data_valid  ;

  output                                          pe21__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane7_strm1_data_mask   ;
  input                                           std__pe21__lane7_strm1_data_valid  ;

  output                                          pe21__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane8_strm0_data_mask   ;
  input                                           std__pe21__lane8_strm0_data_valid  ;

  output                                          pe21__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane8_strm1_data_mask   ;
  input                                           std__pe21__lane8_strm1_data_valid  ;

  output                                          pe21__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane9_strm0_data_mask   ;
  input                                           std__pe21__lane9_strm0_data_valid  ;

  output                                          pe21__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane9_strm1_data_mask   ;
  input                                           std__pe21__lane9_strm1_data_valid  ;

  output                                          pe21__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane10_strm0_data_mask   ;
  input                                           std__pe21__lane10_strm0_data_valid  ;

  output                                          pe21__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane10_strm1_data_mask   ;
  input                                           std__pe21__lane10_strm1_data_valid  ;

  output                                          pe21__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane11_strm0_data_mask   ;
  input                                           std__pe21__lane11_strm0_data_valid  ;

  output                                          pe21__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane11_strm1_data_mask   ;
  input                                           std__pe21__lane11_strm1_data_valid  ;

  output                                          pe21__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane12_strm0_data_mask   ;
  input                                           std__pe21__lane12_strm0_data_valid  ;

  output                                          pe21__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane12_strm1_data_mask   ;
  input                                           std__pe21__lane12_strm1_data_valid  ;

  output                                          pe21__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane13_strm0_data_mask   ;
  input                                           std__pe21__lane13_strm0_data_valid  ;

  output                                          pe21__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane13_strm1_data_mask   ;
  input                                           std__pe21__lane13_strm1_data_valid  ;

  output                                          pe21__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane14_strm0_data_mask   ;
  input                                           std__pe21__lane14_strm0_data_valid  ;

  output                                          pe21__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane14_strm1_data_mask   ;
  input                                           std__pe21__lane14_strm1_data_valid  ;

  output                                          pe21__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane15_strm0_data_mask   ;
  input                                           std__pe21__lane15_strm0_data_valid  ;

  output                                          pe21__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane15_strm1_data_mask   ;
  input                                           std__pe21__lane15_strm1_data_valid  ;

  output                                          pe21__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane16_strm0_data_mask   ;
  input                                           std__pe21__lane16_strm0_data_valid  ;

  output                                          pe21__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane16_strm1_data_mask   ;
  input                                           std__pe21__lane16_strm1_data_valid  ;

  output                                          pe21__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane17_strm0_data_mask   ;
  input                                           std__pe21__lane17_strm0_data_valid  ;

  output                                          pe21__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane17_strm1_data_mask   ;
  input                                           std__pe21__lane17_strm1_data_valid  ;

  output                                          pe21__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane18_strm0_data_mask   ;
  input                                           std__pe21__lane18_strm0_data_valid  ;

  output                                          pe21__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane18_strm1_data_mask   ;
  input                                           std__pe21__lane18_strm1_data_valid  ;

  output                                          pe21__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane19_strm0_data_mask   ;
  input                                           std__pe21__lane19_strm0_data_valid  ;

  output                                          pe21__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane19_strm1_data_mask   ;
  input                                           std__pe21__lane19_strm1_data_valid  ;

  output                                          pe21__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane20_strm0_data_mask   ;
  input                                           std__pe21__lane20_strm0_data_valid  ;

  output                                          pe21__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane20_strm1_data_mask   ;
  input                                           std__pe21__lane20_strm1_data_valid  ;

  output                                          pe21__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane21_strm0_data_mask   ;
  input                                           std__pe21__lane21_strm0_data_valid  ;

  output                                          pe21__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane21_strm1_data_mask   ;
  input                                           std__pe21__lane21_strm1_data_valid  ;

  output                                          pe21__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane22_strm0_data_mask   ;
  input                                           std__pe21__lane22_strm0_data_valid  ;

  output                                          pe21__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane22_strm1_data_mask   ;
  input                                           std__pe21__lane22_strm1_data_valid  ;

  output                                          pe21__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane23_strm0_data_mask   ;
  input                                           std__pe21__lane23_strm0_data_valid  ;

  output                                          pe21__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane23_strm1_data_mask   ;
  input                                           std__pe21__lane23_strm1_data_valid  ;

  output                                          pe21__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane24_strm0_data_mask   ;
  input                                           std__pe21__lane24_strm0_data_valid  ;

  output                                          pe21__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane24_strm1_data_mask   ;
  input                                           std__pe21__lane24_strm1_data_valid  ;

  output                                          pe21__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane25_strm0_data_mask   ;
  input                                           std__pe21__lane25_strm0_data_valid  ;

  output                                          pe21__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane25_strm1_data_mask   ;
  input                                           std__pe21__lane25_strm1_data_valid  ;

  output                                          pe21__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane26_strm0_data_mask   ;
  input                                           std__pe21__lane26_strm0_data_valid  ;

  output                                          pe21__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane26_strm1_data_mask   ;
  input                                           std__pe21__lane26_strm1_data_valid  ;

  output                                          pe21__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane27_strm0_data_mask   ;
  input                                           std__pe21__lane27_strm0_data_valid  ;

  output                                          pe21__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane27_strm1_data_mask   ;
  input                                           std__pe21__lane27_strm1_data_valid  ;

  output                                          pe21__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane28_strm0_data_mask   ;
  input                                           std__pe21__lane28_strm0_data_valid  ;

  output                                          pe21__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane28_strm1_data_mask   ;
  input                                           std__pe21__lane28_strm1_data_valid  ;

  output                                          pe21__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane29_strm0_data_mask   ;
  input                                           std__pe21__lane29_strm0_data_valid  ;

  output                                          pe21__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane29_strm1_data_mask   ;
  input                                           std__pe21__lane29_strm1_data_valid  ;

  output                                          pe21__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane30_strm0_data_mask   ;
  input                                           std__pe21__lane30_strm0_data_valid  ;

  output                                          pe21__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane30_strm1_data_mask   ;
  input                                           std__pe21__lane30_strm1_data_valid  ;

  output                                          pe21__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane31_strm0_data_mask   ;
  input                                           std__pe21__lane31_strm0_data_valid  ;

  output                                          pe21__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe21__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe21__lane31_strm1_data_mask   ;
  input                                           std__pe21__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe22__peId                ;
  input                                         sys__pe22__allSynchronized     ;
  output                                        pe22__sys__thisSynchronized    ;
  output                                        pe22__sys__ready               ;
  output                                        pe22__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe22__oob_cntl            ;
  input                                         std__pe22__oob_valid           ;
  output                                        pe22__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe22__oob_type            ;
  output                                          pe22__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane0_strm0_data_mask   ;
  input                                           std__pe22__lane0_strm0_data_valid  ;

  output                                          pe22__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane0_strm1_data_mask   ;
  input                                           std__pe22__lane0_strm1_data_valid  ;

  output                                          pe22__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane1_strm0_data_mask   ;
  input                                           std__pe22__lane1_strm0_data_valid  ;

  output                                          pe22__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane1_strm1_data_mask   ;
  input                                           std__pe22__lane1_strm1_data_valid  ;

  output                                          pe22__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane2_strm0_data_mask   ;
  input                                           std__pe22__lane2_strm0_data_valid  ;

  output                                          pe22__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane2_strm1_data_mask   ;
  input                                           std__pe22__lane2_strm1_data_valid  ;

  output                                          pe22__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane3_strm0_data_mask   ;
  input                                           std__pe22__lane3_strm0_data_valid  ;

  output                                          pe22__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane3_strm1_data_mask   ;
  input                                           std__pe22__lane3_strm1_data_valid  ;

  output                                          pe22__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane4_strm0_data_mask   ;
  input                                           std__pe22__lane4_strm0_data_valid  ;

  output                                          pe22__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane4_strm1_data_mask   ;
  input                                           std__pe22__lane4_strm1_data_valid  ;

  output                                          pe22__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane5_strm0_data_mask   ;
  input                                           std__pe22__lane5_strm0_data_valid  ;

  output                                          pe22__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane5_strm1_data_mask   ;
  input                                           std__pe22__lane5_strm1_data_valid  ;

  output                                          pe22__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane6_strm0_data_mask   ;
  input                                           std__pe22__lane6_strm0_data_valid  ;

  output                                          pe22__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane6_strm1_data_mask   ;
  input                                           std__pe22__lane6_strm1_data_valid  ;

  output                                          pe22__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane7_strm0_data_mask   ;
  input                                           std__pe22__lane7_strm0_data_valid  ;

  output                                          pe22__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane7_strm1_data_mask   ;
  input                                           std__pe22__lane7_strm1_data_valid  ;

  output                                          pe22__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane8_strm0_data_mask   ;
  input                                           std__pe22__lane8_strm0_data_valid  ;

  output                                          pe22__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane8_strm1_data_mask   ;
  input                                           std__pe22__lane8_strm1_data_valid  ;

  output                                          pe22__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane9_strm0_data_mask   ;
  input                                           std__pe22__lane9_strm0_data_valid  ;

  output                                          pe22__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane9_strm1_data_mask   ;
  input                                           std__pe22__lane9_strm1_data_valid  ;

  output                                          pe22__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane10_strm0_data_mask   ;
  input                                           std__pe22__lane10_strm0_data_valid  ;

  output                                          pe22__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane10_strm1_data_mask   ;
  input                                           std__pe22__lane10_strm1_data_valid  ;

  output                                          pe22__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane11_strm0_data_mask   ;
  input                                           std__pe22__lane11_strm0_data_valid  ;

  output                                          pe22__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane11_strm1_data_mask   ;
  input                                           std__pe22__lane11_strm1_data_valid  ;

  output                                          pe22__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane12_strm0_data_mask   ;
  input                                           std__pe22__lane12_strm0_data_valid  ;

  output                                          pe22__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane12_strm1_data_mask   ;
  input                                           std__pe22__lane12_strm1_data_valid  ;

  output                                          pe22__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane13_strm0_data_mask   ;
  input                                           std__pe22__lane13_strm0_data_valid  ;

  output                                          pe22__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane13_strm1_data_mask   ;
  input                                           std__pe22__lane13_strm1_data_valid  ;

  output                                          pe22__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane14_strm0_data_mask   ;
  input                                           std__pe22__lane14_strm0_data_valid  ;

  output                                          pe22__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane14_strm1_data_mask   ;
  input                                           std__pe22__lane14_strm1_data_valid  ;

  output                                          pe22__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane15_strm0_data_mask   ;
  input                                           std__pe22__lane15_strm0_data_valid  ;

  output                                          pe22__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane15_strm1_data_mask   ;
  input                                           std__pe22__lane15_strm1_data_valid  ;

  output                                          pe22__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane16_strm0_data_mask   ;
  input                                           std__pe22__lane16_strm0_data_valid  ;

  output                                          pe22__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane16_strm1_data_mask   ;
  input                                           std__pe22__lane16_strm1_data_valid  ;

  output                                          pe22__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane17_strm0_data_mask   ;
  input                                           std__pe22__lane17_strm0_data_valid  ;

  output                                          pe22__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane17_strm1_data_mask   ;
  input                                           std__pe22__lane17_strm1_data_valid  ;

  output                                          pe22__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane18_strm0_data_mask   ;
  input                                           std__pe22__lane18_strm0_data_valid  ;

  output                                          pe22__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane18_strm1_data_mask   ;
  input                                           std__pe22__lane18_strm1_data_valid  ;

  output                                          pe22__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane19_strm0_data_mask   ;
  input                                           std__pe22__lane19_strm0_data_valid  ;

  output                                          pe22__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane19_strm1_data_mask   ;
  input                                           std__pe22__lane19_strm1_data_valid  ;

  output                                          pe22__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane20_strm0_data_mask   ;
  input                                           std__pe22__lane20_strm0_data_valid  ;

  output                                          pe22__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane20_strm1_data_mask   ;
  input                                           std__pe22__lane20_strm1_data_valid  ;

  output                                          pe22__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane21_strm0_data_mask   ;
  input                                           std__pe22__lane21_strm0_data_valid  ;

  output                                          pe22__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane21_strm1_data_mask   ;
  input                                           std__pe22__lane21_strm1_data_valid  ;

  output                                          pe22__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane22_strm0_data_mask   ;
  input                                           std__pe22__lane22_strm0_data_valid  ;

  output                                          pe22__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane22_strm1_data_mask   ;
  input                                           std__pe22__lane22_strm1_data_valid  ;

  output                                          pe22__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane23_strm0_data_mask   ;
  input                                           std__pe22__lane23_strm0_data_valid  ;

  output                                          pe22__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane23_strm1_data_mask   ;
  input                                           std__pe22__lane23_strm1_data_valid  ;

  output                                          pe22__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane24_strm0_data_mask   ;
  input                                           std__pe22__lane24_strm0_data_valid  ;

  output                                          pe22__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane24_strm1_data_mask   ;
  input                                           std__pe22__lane24_strm1_data_valid  ;

  output                                          pe22__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane25_strm0_data_mask   ;
  input                                           std__pe22__lane25_strm0_data_valid  ;

  output                                          pe22__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane25_strm1_data_mask   ;
  input                                           std__pe22__lane25_strm1_data_valid  ;

  output                                          pe22__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane26_strm0_data_mask   ;
  input                                           std__pe22__lane26_strm0_data_valid  ;

  output                                          pe22__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane26_strm1_data_mask   ;
  input                                           std__pe22__lane26_strm1_data_valid  ;

  output                                          pe22__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane27_strm0_data_mask   ;
  input                                           std__pe22__lane27_strm0_data_valid  ;

  output                                          pe22__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane27_strm1_data_mask   ;
  input                                           std__pe22__lane27_strm1_data_valid  ;

  output                                          pe22__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane28_strm0_data_mask   ;
  input                                           std__pe22__lane28_strm0_data_valid  ;

  output                                          pe22__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane28_strm1_data_mask   ;
  input                                           std__pe22__lane28_strm1_data_valid  ;

  output                                          pe22__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane29_strm0_data_mask   ;
  input                                           std__pe22__lane29_strm0_data_valid  ;

  output                                          pe22__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane29_strm1_data_mask   ;
  input                                           std__pe22__lane29_strm1_data_valid  ;

  output                                          pe22__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane30_strm0_data_mask   ;
  input                                           std__pe22__lane30_strm0_data_valid  ;

  output                                          pe22__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane30_strm1_data_mask   ;
  input                                           std__pe22__lane30_strm1_data_valid  ;

  output                                          pe22__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane31_strm0_data_mask   ;
  input                                           std__pe22__lane31_strm0_data_valid  ;

  output                                          pe22__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe22__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe22__lane31_strm1_data_mask   ;
  input                                           std__pe22__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe23__peId                ;
  input                                         sys__pe23__allSynchronized     ;
  output                                        pe23__sys__thisSynchronized    ;
  output                                        pe23__sys__ready               ;
  output                                        pe23__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe23__oob_cntl            ;
  input                                         std__pe23__oob_valid           ;
  output                                        pe23__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe23__oob_type            ;
  output                                          pe23__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane0_strm0_data_mask   ;
  input                                           std__pe23__lane0_strm0_data_valid  ;

  output                                          pe23__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane0_strm1_data_mask   ;
  input                                           std__pe23__lane0_strm1_data_valid  ;

  output                                          pe23__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane1_strm0_data_mask   ;
  input                                           std__pe23__lane1_strm0_data_valid  ;

  output                                          pe23__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane1_strm1_data_mask   ;
  input                                           std__pe23__lane1_strm1_data_valid  ;

  output                                          pe23__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane2_strm0_data_mask   ;
  input                                           std__pe23__lane2_strm0_data_valid  ;

  output                                          pe23__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane2_strm1_data_mask   ;
  input                                           std__pe23__lane2_strm1_data_valid  ;

  output                                          pe23__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane3_strm0_data_mask   ;
  input                                           std__pe23__lane3_strm0_data_valid  ;

  output                                          pe23__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane3_strm1_data_mask   ;
  input                                           std__pe23__lane3_strm1_data_valid  ;

  output                                          pe23__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane4_strm0_data_mask   ;
  input                                           std__pe23__lane4_strm0_data_valid  ;

  output                                          pe23__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane4_strm1_data_mask   ;
  input                                           std__pe23__lane4_strm1_data_valid  ;

  output                                          pe23__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane5_strm0_data_mask   ;
  input                                           std__pe23__lane5_strm0_data_valid  ;

  output                                          pe23__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane5_strm1_data_mask   ;
  input                                           std__pe23__lane5_strm1_data_valid  ;

  output                                          pe23__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane6_strm0_data_mask   ;
  input                                           std__pe23__lane6_strm0_data_valid  ;

  output                                          pe23__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane6_strm1_data_mask   ;
  input                                           std__pe23__lane6_strm1_data_valid  ;

  output                                          pe23__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane7_strm0_data_mask   ;
  input                                           std__pe23__lane7_strm0_data_valid  ;

  output                                          pe23__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane7_strm1_data_mask   ;
  input                                           std__pe23__lane7_strm1_data_valid  ;

  output                                          pe23__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane8_strm0_data_mask   ;
  input                                           std__pe23__lane8_strm0_data_valid  ;

  output                                          pe23__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane8_strm1_data_mask   ;
  input                                           std__pe23__lane8_strm1_data_valid  ;

  output                                          pe23__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane9_strm0_data_mask   ;
  input                                           std__pe23__lane9_strm0_data_valid  ;

  output                                          pe23__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane9_strm1_data_mask   ;
  input                                           std__pe23__lane9_strm1_data_valid  ;

  output                                          pe23__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane10_strm0_data_mask   ;
  input                                           std__pe23__lane10_strm0_data_valid  ;

  output                                          pe23__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane10_strm1_data_mask   ;
  input                                           std__pe23__lane10_strm1_data_valid  ;

  output                                          pe23__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane11_strm0_data_mask   ;
  input                                           std__pe23__lane11_strm0_data_valid  ;

  output                                          pe23__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane11_strm1_data_mask   ;
  input                                           std__pe23__lane11_strm1_data_valid  ;

  output                                          pe23__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane12_strm0_data_mask   ;
  input                                           std__pe23__lane12_strm0_data_valid  ;

  output                                          pe23__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane12_strm1_data_mask   ;
  input                                           std__pe23__lane12_strm1_data_valid  ;

  output                                          pe23__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane13_strm0_data_mask   ;
  input                                           std__pe23__lane13_strm0_data_valid  ;

  output                                          pe23__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane13_strm1_data_mask   ;
  input                                           std__pe23__lane13_strm1_data_valid  ;

  output                                          pe23__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane14_strm0_data_mask   ;
  input                                           std__pe23__lane14_strm0_data_valid  ;

  output                                          pe23__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane14_strm1_data_mask   ;
  input                                           std__pe23__lane14_strm1_data_valid  ;

  output                                          pe23__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane15_strm0_data_mask   ;
  input                                           std__pe23__lane15_strm0_data_valid  ;

  output                                          pe23__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane15_strm1_data_mask   ;
  input                                           std__pe23__lane15_strm1_data_valid  ;

  output                                          pe23__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane16_strm0_data_mask   ;
  input                                           std__pe23__lane16_strm0_data_valid  ;

  output                                          pe23__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane16_strm1_data_mask   ;
  input                                           std__pe23__lane16_strm1_data_valid  ;

  output                                          pe23__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane17_strm0_data_mask   ;
  input                                           std__pe23__lane17_strm0_data_valid  ;

  output                                          pe23__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane17_strm1_data_mask   ;
  input                                           std__pe23__lane17_strm1_data_valid  ;

  output                                          pe23__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane18_strm0_data_mask   ;
  input                                           std__pe23__lane18_strm0_data_valid  ;

  output                                          pe23__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane18_strm1_data_mask   ;
  input                                           std__pe23__lane18_strm1_data_valid  ;

  output                                          pe23__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane19_strm0_data_mask   ;
  input                                           std__pe23__lane19_strm0_data_valid  ;

  output                                          pe23__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane19_strm1_data_mask   ;
  input                                           std__pe23__lane19_strm1_data_valid  ;

  output                                          pe23__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane20_strm0_data_mask   ;
  input                                           std__pe23__lane20_strm0_data_valid  ;

  output                                          pe23__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane20_strm1_data_mask   ;
  input                                           std__pe23__lane20_strm1_data_valid  ;

  output                                          pe23__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane21_strm0_data_mask   ;
  input                                           std__pe23__lane21_strm0_data_valid  ;

  output                                          pe23__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane21_strm1_data_mask   ;
  input                                           std__pe23__lane21_strm1_data_valid  ;

  output                                          pe23__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane22_strm0_data_mask   ;
  input                                           std__pe23__lane22_strm0_data_valid  ;

  output                                          pe23__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane22_strm1_data_mask   ;
  input                                           std__pe23__lane22_strm1_data_valid  ;

  output                                          pe23__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane23_strm0_data_mask   ;
  input                                           std__pe23__lane23_strm0_data_valid  ;

  output                                          pe23__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane23_strm1_data_mask   ;
  input                                           std__pe23__lane23_strm1_data_valid  ;

  output                                          pe23__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane24_strm0_data_mask   ;
  input                                           std__pe23__lane24_strm0_data_valid  ;

  output                                          pe23__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane24_strm1_data_mask   ;
  input                                           std__pe23__lane24_strm1_data_valid  ;

  output                                          pe23__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane25_strm0_data_mask   ;
  input                                           std__pe23__lane25_strm0_data_valid  ;

  output                                          pe23__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane25_strm1_data_mask   ;
  input                                           std__pe23__lane25_strm1_data_valid  ;

  output                                          pe23__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane26_strm0_data_mask   ;
  input                                           std__pe23__lane26_strm0_data_valid  ;

  output                                          pe23__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane26_strm1_data_mask   ;
  input                                           std__pe23__lane26_strm1_data_valid  ;

  output                                          pe23__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane27_strm0_data_mask   ;
  input                                           std__pe23__lane27_strm0_data_valid  ;

  output                                          pe23__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane27_strm1_data_mask   ;
  input                                           std__pe23__lane27_strm1_data_valid  ;

  output                                          pe23__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane28_strm0_data_mask   ;
  input                                           std__pe23__lane28_strm0_data_valid  ;

  output                                          pe23__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane28_strm1_data_mask   ;
  input                                           std__pe23__lane28_strm1_data_valid  ;

  output                                          pe23__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane29_strm0_data_mask   ;
  input                                           std__pe23__lane29_strm0_data_valid  ;

  output                                          pe23__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane29_strm1_data_mask   ;
  input                                           std__pe23__lane29_strm1_data_valid  ;

  output                                          pe23__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane30_strm0_data_mask   ;
  input                                           std__pe23__lane30_strm0_data_valid  ;

  output                                          pe23__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane30_strm1_data_mask   ;
  input                                           std__pe23__lane30_strm1_data_valid  ;

  output                                          pe23__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane31_strm0_data_mask   ;
  input                                           std__pe23__lane31_strm0_data_valid  ;

  output                                          pe23__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe23__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe23__lane31_strm1_data_mask   ;
  input                                           std__pe23__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe24__peId                ;
  input                                         sys__pe24__allSynchronized     ;
  output                                        pe24__sys__thisSynchronized    ;
  output                                        pe24__sys__ready               ;
  output                                        pe24__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe24__oob_cntl            ;
  input                                         std__pe24__oob_valid           ;
  output                                        pe24__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe24__oob_type            ;
  output                                          pe24__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane0_strm0_data_mask   ;
  input                                           std__pe24__lane0_strm0_data_valid  ;

  output                                          pe24__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane0_strm1_data_mask   ;
  input                                           std__pe24__lane0_strm1_data_valid  ;

  output                                          pe24__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane1_strm0_data_mask   ;
  input                                           std__pe24__lane1_strm0_data_valid  ;

  output                                          pe24__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane1_strm1_data_mask   ;
  input                                           std__pe24__lane1_strm1_data_valid  ;

  output                                          pe24__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane2_strm0_data_mask   ;
  input                                           std__pe24__lane2_strm0_data_valid  ;

  output                                          pe24__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane2_strm1_data_mask   ;
  input                                           std__pe24__lane2_strm1_data_valid  ;

  output                                          pe24__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane3_strm0_data_mask   ;
  input                                           std__pe24__lane3_strm0_data_valid  ;

  output                                          pe24__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane3_strm1_data_mask   ;
  input                                           std__pe24__lane3_strm1_data_valid  ;

  output                                          pe24__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane4_strm0_data_mask   ;
  input                                           std__pe24__lane4_strm0_data_valid  ;

  output                                          pe24__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane4_strm1_data_mask   ;
  input                                           std__pe24__lane4_strm1_data_valid  ;

  output                                          pe24__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane5_strm0_data_mask   ;
  input                                           std__pe24__lane5_strm0_data_valid  ;

  output                                          pe24__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane5_strm1_data_mask   ;
  input                                           std__pe24__lane5_strm1_data_valid  ;

  output                                          pe24__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane6_strm0_data_mask   ;
  input                                           std__pe24__lane6_strm0_data_valid  ;

  output                                          pe24__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane6_strm1_data_mask   ;
  input                                           std__pe24__lane6_strm1_data_valid  ;

  output                                          pe24__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane7_strm0_data_mask   ;
  input                                           std__pe24__lane7_strm0_data_valid  ;

  output                                          pe24__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane7_strm1_data_mask   ;
  input                                           std__pe24__lane7_strm1_data_valid  ;

  output                                          pe24__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane8_strm0_data_mask   ;
  input                                           std__pe24__lane8_strm0_data_valid  ;

  output                                          pe24__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane8_strm1_data_mask   ;
  input                                           std__pe24__lane8_strm1_data_valid  ;

  output                                          pe24__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane9_strm0_data_mask   ;
  input                                           std__pe24__lane9_strm0_data_valid  ;

  output                                          pe24__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane9_strm1_data_mask   ;
  input                                           std__pe24__lane9_strm1_data_valid  ;

  output                                          pe24__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane10_strm0_data_mask   ;
  input                                           std__pe24__lane10_strm0_data_valid  ;

  output                                          pe24__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane10_strm1_data_mask   ;
  input                                           std__pe24__lane10_strm1_data_valid  ;

  output                                          pe24__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane11_strm0_data_mask   ;
  input                                           std__pe24__lane11_strm0_data_valid  ;

  output                                          pe24__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane11_strm1_data_mask   ;
  input                                           std__pe24__lane11_strm1_data_valid  ;

  output                                          pe24__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane12_strm0_data_mask   ;
  input                                           std__pe24__lane12_strm0_data_valid  ;

  output                                          pe24__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane12_strm1_data_mask   ;
  input                                           std__pe24__lane12_strm1_data_valid  ;

  output                                          pe24__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane13_strm0_data_mask   ;
  input                                           std__pe24__lane13_strm0_data_valid  ;

  output                                          pe24__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane13_strm1_data_mask   ;
  input                                           std__pe24__lane13_strm1_data_valid  ;

  output                                          pe24__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane14_strm0_data_mask   ;
  input                                           std__pe24__lane14_strm0_data_valid  ;

  output                                          pe24__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane14_strm1_data_mask   ;
  input                                           std__pe24__lane14_strm1_data_valid  ;

  output                                          pe24__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane15_strm0_data_mask   ;
  input                                           std__pe24__lane15_strm0_data_valid  ;

  output                                          pe24__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane15_strm1_data_mask   ;
  input                                           std__pe24__lane15_strm1_data_valid  ;

  output                                          pe24__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane16_strm0_data_mask   ;
  input                                           std__pe24__lane16_strm0_data_valid  ;

  output                                          pe24__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane16_strm1_data_mask   ;
  input                                           std__pe24__lane16_strm1_data_valid  ;

  output                                          pe24__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane17_strm0_data_mask   ;
  input                                           std__pe24__lane17_strm0_data_valid  ;

  output                                          pe24__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane17_strm1_data_mask   ;
  input                                           std__pe24__lane17_strm1_data_valid  ;

  output                                          pe24__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane18_strm0_data_mask   ;
  input                                           std__pe24__lane18_strm0_data_valid  ;

  output                                          pe24__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane18_strm1_data_mask   ;
  input                                           std__pe24__lane18_strm1_data_valid  ;

  output                                          pe24__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane19_strm0_data_mask   ;
  input                                           std__pe24__lane19_strm0_data_valid  ;

  output                                          pe24__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane19_strm1_data_mask   ;
  input                                           std__pe24__lane19_strm1_data_valid  ;

  output                                          pe24__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane20_strm0_data_mask   ;
  input                                           std__pe24__lane20_strm0_data_valid  ;

  output                                          pe24__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane20_strm1_data_mask   ;
  input                                           std__pe24__lane20_strm1_data_valid  ;

  output                                          pe24__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane21_strm0_data_mask   ;
  input                                           std__pe24__lane21_strm0_data_valid  ;

  output                                          pe24__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane21_strm1_data_mask   ;
  input                                           std__pe24__lane21_strm1_data_valid  ;

  output                                          pe24__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane22_strm0_data_mask   ;
  input                                           std__pe24__lane22_strm0_data_valid  ;

  output                                          pe24__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane22_strm1_data_mask   ;
  input                                           std__pe24__lane22_strm1_data_valid  ;

  output                                          pe24__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane23_strm0_data_mask   ;
  input                                           std__pe24__lane23_strm0_data_valid  ;

  output                                          pe24__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane23_strm1_data_mask   ;
  input                                           std__pe24__lane23_strm1_data_valid  ;

  output                                          pe24__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane24_strm0_data_mask   ;
  input                                           std__pe24__lane24_strm0_data_valid  ;

  output                                          pe24__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane24_strm1_data_mask   ;
  input                                           std__pe24__lane24_strm1_data_valid  ;

  output                                          pe24__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane25_strm0_data_mask   ;
  input                                           std__pe24__lane25_strm0_data_valid  ;

  output                                          pe24__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane25_strm1_data_mask   ;
  input                                           std__pe24__lane25_strm1_data_valid  ;

  output                                          pe24__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane26_strm0_data_mask   ;
  input                                           std__pe24__lane26_strm0_data_valid  ;

  output                                          pe24__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane26_strm1_data_mask   ;
  input                                           std__pe24__lane26_strm1_data_valid  ;

  output                                          pe24__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane27_strm0_data_mask   ;
  input                                           std__pe24__lane27_strm0_data_valid  ;

  output                                          pe24__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane27_strm1_data_mask   ;
  input                                           std__pe24__lane27_strm1_data_valid  ;

  output                                          pe24__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane28_strm0_data_mask   ;
  input                                           std__pe24__lane28_strm0_data_valid  ;

  output                                          pe24__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane28_strm1_data_mask   ;
  input                                           std__pe24__lane28_strm1_data_valid  ;

  output                                          pe24__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane29_strm0_data_mask   ;
  input                                           std__pe24__lane29_strm0_data_valid  ;

  output                                          pe24__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane29_strm1_data_mask   ;
  input                                           std__pe24__lane29_strm1_data_valid  ;

  output                                          pe24__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane30_strm0_data_mask   ;
  input                                           std__pe24__lane30_strm0_data_valid  ;

  output                                          pe24__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane30_strm1_data_mask   ;
  input                                           std__pe24__lane30_strm1_data_valid  ;

  output                                          pe24__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane31_strm0_data_mask   ;
  input                                           std__pe24__lane31_strm0_data_valid  ;

  output                                          pe24__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe24__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe24__lane31_strm1_data_mask   ;
  input                                           std__pe24__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe25__peId                ;
  input                                         sys__pe25__allSynchronized     ;
  output                                        pe25__sys__thisSynchronized    ;
  output                                        pe25__sys__ready               ;
  output                                        pe25__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe25__oob_cntl            ;
  input                                         std__pe25__oob_valid           ;
  output                                        pe25__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe25__oob_type            ;
  output                                          pe25__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane0_strm0_data_mask   ;
  input                                           std__pe25__lane0_strm0_data_valid  ;

  output                                          pe25__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane0_strm1_data_mask   ;
  input                                           std__pe25__lane0_strm1_data_valid  ;

  output                                          pe25__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane1_strm0_data_mask   ;
  input                                           std__pe25__lane1_strm0_data_valid  ;

  output                                          pe25__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane1_strm1_data_mask   ;
  input                                           std__pe25__lane1_strm1_data_valid  ;

  output                                          pe25__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane2_strm0_data_mask   ;
  input                                           std__pe25__lane2_strm0_data_valid  ;

  output                                          pe25__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane2_strm1_data_mask   ;
  input                                           std__pe25__lane2_strm1_data_valid  ;

  output                                          pe25__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane3_strm0_data_mask   ;
  input                                           std__pe25__lane3_strm0_data_valid  ;

  output                                          pe25__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane3_strm1_data_mask   ;
  input                                           std__pe25__lane3_strm1_data_valid  ;

  output                                          pe25__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane4_strm0_data_mask   ;
  input                                           std__pe25__lane4_strm0_data_valid  ;

  output                                          pe25__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane4_strm1_data_mask   ;
  input                                           std__pe25__lane4_strm1_data_valid  ;

  output                                          pe25__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane5_strm0_data_mask   ;
  input                                           std__pe25__lane5_strm0_data_valid  ;

  output                                          pe25__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane5_strm1_data_mask   ;
  input                                           std__pe25__lane5_strm1_data_valid  ;

  output                                          pe25__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane6_strm0_data_mask   ;
  input                                           std__pe25__lane6_strm0_data_valid  ;

  output                                          pe25__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane6_strm1_data_mask   ;
  input                                           std__pe25__lane6_strm1_data_valid  ;

  output                                          pe25__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane7_strm0_data_mask   ;
  input                                           std__pe25__lane7_strm0_data_valid  ;

  output                                          pe25__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane7_strm1_data_mask   ;
  input                                           std__pe25__lane7_strm1_data_valid  ;

  output                                          pe25__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane8_strm0_data_mask   ;
  input                                           std__pe25__lane8_strm0_data_valid  ;

  output                                          pe25__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane8_strm1_data_mask   ;
  input                                           std__pe25__lane8_strm1_data_valid  ;

  output                                          pe25__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane9_strm0_data_mask   ;
  input                                           std__pe25__lane9_strm0_data_valid  ;

  output                                          pe25__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane9_strm1_data_mask   ;
  input                                           std__pe25__lane9_strm1_data_valid  ;

  output                                          pe25__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane10_strm0_data_mask   ;
  input                                           std__pe25__lane10_strm0_data_valid  ;

  output                                          pe25__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane10_strm1_data_mask   ;
  input                                           std__pe25__lane10_strm1_data_valid  ;

  output                                          pe25__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane11_strm0_data_mask   ;
  input                                           std__pe25__lane11_strm0_data_valid  ;

  output                                          pe25__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane11_strm1_data_mask   ;
  input                                           std__pe25__lane11_strm1_data_valid  ;

  output                                          pe25__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane12_strm0_data_mask   ;
  input                                           std__pe25__lane12_strm0_data_valid  ;

  output                                          pe25__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane12_strm1_data_mask   ;
  input                                           std__pe25__lane12_strm1_data_valid  ;

  output                                          pe25__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane13_strm0_data_mask   ;
  input                                           std__pe25__lane13_strm0_data_valid  ;

  output                                          pe25__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane13_strm1_data_mask   ;
  input                                           std__pe25__lane13_strm1_data_valid  ;

  output                                          pe25__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane14_strm0_data_mask   ;
  input                                           std__pe25__lane14_strm0_data_valid  ;

  output                                          pe25__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane14_strm1_data_mask   ;
  input                                           std__pe25__lane14_strm1_data_valid  ;

  output                                          pe25__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane15_strm0_data_mask   ;
  input                                           std__pe25__lane15_strm0_data_valid  ;

  output                                          pe25__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane15_strm1_data_mask   ;
  input                                           std__pe25__lane15_strm1_data_valid  ;

  output                                          pe25__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane16_strm0_data_mask   ;
  input                                           std__pe25__lane16_strm0_data_valid  ;

  output                                          pe25__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane16_strm1_data_mask   ;
  input                                           std__pe25__lane16_strm1_data_valid  ;

  output                                          pe25__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane17_strm0_data_mask   ;
  input                                           std__pe25__lane17_strm0_data_valid  ;

  output                                          pe25__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane17_strm1_data_mask   ;
  input                                           std__pe25__lane17_strm1_data_valid  ;

  output                                          pe25__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane18_strm0_data_mask   ;
  input                                           std__pe25__lane18_strm0_data_valid  ;

  output                                          pe25__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane18_strm1_data_mask   ;
  input                                           std__pe25__lane18_strm1_data_valid  ;

  output                                          pe25__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane19_strm0_data_mask   ;
  input                                           std__pe25__lane19_strm0_data_valid  ;

  output                                          pe25__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane19_strm1_data_mask   ;
  input                                           std__pe25__lane19_strm1_data_valid  ;

  output                                          pe25__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane20_strm0_data_mask   ;
  input                                           std__pe25__lane20_strm0_data_valid  ;

  output                                          pe25__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane20_strm1_data_mask   ;
  input                                           std__pe25__lane20_strm1_data_valid  ;

  output                                          pe25__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane21_strm0_data_mask   ;
  input                                           std__pe25__lane21_strm0_data_valid  ;

  output                                          pe25__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane21_strm1_data_mask   ;
  input                                           std__pe25__lane21_strm1_data_valid  ;

  output                                          pe25__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane22_strm0_data_mask   ;
  input                                           std__pe25__lane22_strm0_data_valid  ;

  output                                          pe25__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane22_strm1_data_mask   ;
  input                                           std__pe25__lane22_strm1_data_valid  ;

  output                                          pe25__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane23_strm0_data_mask   ;
  input                                           std__pe25__lane23_strm0_data_valid  ;

  output                                          pe25__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane23_strm1_data_mask   ;
  input                                           std__pe25__lane23_strm1_data_valid  ;

  output                                          pe25__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane24_strm0_data_mask   ;
  input                                           std__pe25__lane24_strm0_data_valid  ;

  output                                          pe25__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane24_strm1_data_mask   ;
  input                                           std__pe25__lane24_strm1_data_valid  ;

  output                                          pe25__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane25_strm0_data_mask   ;
  input                                           std__pe25__lane25_strm0_data_valid  ;

  output                                          pe25__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane25_strm1_data_mask   ;
  input                                           std__pe25__lane25_strm1_data_valid  ;

  output                                          pe25__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane26_strm0_data_mask   ;
  input                                           std__pe25__lane26_strm0_data_valid  ;

  output                                          pe25__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane26_strm1_data_mask   ;
  input                                           std__pe25__lane26_strm1_data_valid  ;

  output                                          pe25__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane27_strm0_data_mask   ;
  input                                           std__pe25__lane27_strm0_data_valid  ;

  output                                          pe25__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane27_strm1_data_mask   ;
  input                                           std__pe25__lane27_strm1_data_valid  ;

  output                                          pe25__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane28_strm0_data_mask   ;
  input                                           std__pe25__lane28_strm0_data_valid  ;

  output                                          pe25__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane28_strm1_data_mask   ;
  input                                           std__pe25__lane28_strm1_data_valid  ;

  output                                          pe25__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane29_strm0_data_mask   ;
  input                                           std__pe25__lane29_strm0_data_valid  ;

  output                                          pe25__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane29_strm1_data_mask   ;
  input                                           std__pe25__lane29_strm1_data_valid  ;

  output                                          pe25__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane30_strm0_data_mask   ;
  input                                           std__pe25__lane30_strm0_data_valid  ;

  output                                          pe25__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane30_strm1_data_mask   ;
  input                                           std__pe25__lane30_strm1_data_valid  ;

  output                                          pe25__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane31_strm0_data_mask   ;
  input                                           std__pe25__lane31_strm0_data_valid  ;

  output                                          pe25__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe25__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe25__lane31_strm1_data_mask   ;
  input                                           std__pe25__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe26__peId                ;
  input                                         sys__pe26__allSynchronized     ;
  output                                        pe26__sys__thisSynchronized    ;
  output                                        pe26__sys__ready               ;
  output                                        pe26__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe26__oob_cntl            ;
  input                                         std__pe26__oob_valid           ;
  output                                        pe26__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe26__oob_type            ;
  output                                          pe26__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane0_strm0_data_mask   ;
  input                                           std__pe26__lane0_strm0_data_valid  ;

  output                                          pe26__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane0_strm1_data_mask   ;
  input                                           std__pe26__lane0_strm1_data_valid  ;

  output                                          pe26__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane1_strm0_data_mask   ;
  input                                           std__pe26__lane1_strm0_data_valid  ;

  output                                          pe26__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane1_strm1_data_mask   ;
  input                                           std__pe26__lane1_strm1_data_valid  ;

  output                                          pe26__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane2_strm0_data_mask   ;
  input                                           std__pe26__lane2_strm0_data_valid  ;

  output                                          pe26__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane2_strm1_data_mask   ;
  input                                           std__pe26__lane2_strm1_data_valid  ;

  output                                          pe26__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane3_strm0_data_mask   ;
  input                                           std__pe26__lane3_strm0_data_valid  ;

  output                                          pe26__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane3_strm1_data_mask   ;
  input                                           std__pe26__lane3_strm1_data_valid  ;

  output                                          pe26__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane4_strm0_data_mask   ;
  input                                           std__pe26__lane4_strm0_data_valid  ;

  output                                          pe26__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane4_strm1_data_mask   ;
  input                                           std__pe26__lane4_strm1_data_valid  ;

  output                                          pe26__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane5_strm0_data_mask   ;
  input                                           std__pe26__lane5_strm0_data_valid  ;

  output                                          pe26__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane5_strm1_data_mask   ;
  input                                           std__pe26__lane5_strm1_data_valid  ;

  output                                          pe26__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane6_strm0_data_mask   ;
  input                                           std__pe26__lane6_strm0_data_valid  ;

  output                                          pe26__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane6_strm1_data_mask   ;
  input                                           std__pe26__lane6_strm1_data_valid  ;

  output                                          pe26__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane7_strm0_data_mask   ;
  input                                           std__pe26__lane7_strm0_data_valid  ;

  output                                          pe26__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane7_strm1_data_mask   ;
  input                                           std__pe26__lane7_strm1_data_valid  ;

  output                                          pe26__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane8_strm0_data_mask   ;
  input                                           std__pe26__lane8_strm0_data_valid  ;

  output                                          pe26__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane8_strm1_data_mask   ;
  input                                           std__pe26__lane8_strm1_data_valid  ;

  output                                          pe26__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane9_strm0_data_mask   ;
  input                                           std__pe26__lane9_strm0_data_valid  ;

  output                                          pe26__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane9_strm1_data_mask   ;
  input                                           std__pe26__lane9_strm1_data_valid  ;

  output                                          pe26__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane10_strm0_data_mask   ;
  input                                           std__pe26__lane10_strm0_data_valid  ;

  output                                          pe26__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane10_strm1_data_mask   ;
  input                                           std__pe26__lane10_strm1_data_valid  ;

  output                                          pe26__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane11_strm0_data_mask   ;
  input                                           std__pe26__lane11_strm0_data_valid  ;

  output                                          pe26__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane11_strm1_data_mask   ;
  input                                           std__pe26__lane11_strm1_data_valid  ;

  output                                          pe26__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane12_strm0_data_mask   ;
  input                                           std__pe26__lane12_strm0_data_valid  ;

  output                                          pe26__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane12_strm1_data_mask   ;
  input                                           std__pe26__lane12_strm1_data_valid  ;

  output                                          pe26__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane13_strm0_data_mask   ;
  input                                           std__pe26__lane13_strm0_data_valid  ;

  output                                          pe26__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane13_strm1_data_mask   ;
  input                                           std__pe26__lane13_strm1_data_valid  ;

  output                                          pe26__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane14_strm0_data_mask   ;
  input                                           std__pe26__lane14_strm0_data_valid  ;

  output                                          pe26__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane14_strm1_data_mask   ;
  input                                           std__pe26__lane14_strm1_data_valid  ;

  output                                          pe26__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane15_strm0_data_mask   ;
  input                                           std__pe26__lane15_strm0_data_valid  ;

  output                                          pe26__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane15_strm1_data_mask   ;
  input                                           std__pe26__lane15_strm1_data_valid  ;

  output                                          pe26__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane16_strm0_data_mask   ;
  input                                           std__pe26__lane16_strm0_data_valid  ;

  output                                          pe26__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane16_strm1_data_mask   ;
  input                                           std__pe26__lane16_strm1_data_valid  ;

  output                                          pe26__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane17_strm0_data_mask   ;
  input                                           std__pe26__lane17_strm0_data_valid  ;

  output                                          pe26__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane17_strm1_data_mask   ;
  input                                           std__pe26__lane17_strm1_data_valid  ;

  output                                          pe26__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane18_strm0_data_mask   ;
  input                                           std__pe26__lane18_strm0_data_valid  ;

  output                                          pe26__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane18_strm1_data_mask   ;
  input                                           std__pe26__lane18_strm1_data_valid  ;

  output                                          pe26__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane19_strm0_data_mask   ;
  input                                           std__pe26__lane19_strm0_data_valid  ;

  output                                          pe26__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane19_strm1_data_mask   ;
  input                                           std__pe26__lane19_strm1_data_valid  ;

  output                                          pe26__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane20_strm0_data_mask   ;
  input                                           std__pe26__lane20_strm0_data_valid  ;

  output                                          pe26__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane20_strm1_data_mask   ;
  input                                           std__pe26__lane20_strm1_data_valid  ;

  output                                          pe26__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane21_strm0_data_mask   ;
  input                                           std__pe26__lane21_strm0_data_valid  ;

  output                                          pe26__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane21_strm1_data_mask   ;
  input                                           std__pe26__lane21_strm1_data_valid  ;

  output                                          pe26__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane22_strm0_data_mask   ;
  input                                           std__pe26__lane22_strm0_data_valid  ;

  output                                          pe26__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane22_strm1_data_mask   ;
  input                                           std__pe26__lane22_strm1_data_valid  ;

  output                                          pe26__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane23_strm0_data_mask   ;
  input                                           std__pe26__lane23_strm0_data_valid  ;

  output                                          pe26__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane23_strm1_data_mask   ;
  input                                           std__pe26__lane23_strm1_data_valid  ;

  output                                          pe26__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane24_strm0_data_mask   ;
  input                                           std__pe26__lane24_strm0_data_valid  ;

  output                                          pe26__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane24_strm1_data_mask   ;
  input                                           std__pe26__lane24_strm1_data_valid  ;

  output                                          pe26__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane25_strm0_data_mask   ;
  input                                           std__pe26__lane25_strm0_data_valid  ;

  output                                          pe26__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane25_strm1_data_mask   ;
  input                                           std__pe26__lane25_strm1_data_valid  ;

  output                                          pe26__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane26_strm0_data_mask   ;
  input                                           std__pe26__lane26_strm0_data_valid  ;

  output                                          pe26__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane26_strm1_data_mask   ;
  input                                           std__pe26__lane26_strm1_data_valid  ;

  output                                          pe26__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane27_strm0_data_mask   ;
  input                                           std__pe26__lane27_strm0_data_valid  ;

  output                                          pe26__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane27_strm1_data_mask   ;
  input                                           std__pe26__lane27_strm1_data_valid  ;

  output                                          pe26__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane28_strm0_data_mask   ;
  input                                           std__pe26__lane28_strm0_data_valid  ;

  output                                          pe26__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane28_strm1_data_mask   ;
  input                                           std__pe26__lane28_strm1_data_valid  ;

  output                                          pe26__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane29_strm0_data_mask   ;
  input                                           std__pe26__lane29_strm0_data_valid  ;

  output                                          pe26__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane29_strm1_data_mask   ;
  input                                           std__pe26__lane29_strm1_data_valid  ;

  output                                          pe26__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane30_strm0_data_mask   ;
  input                                           std__pe26__lane30_strm0_data_valid  ;

  output                                          pe26__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane30_strm1_data_mask   ;
  input                                           std__pe26__lane30_strm1_data_valid  ;

  output                                          pe26__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane31_strm0_data_mask   ;
  input                                           std__pe26__lane31_strm0_data_valid  ;

  output                                          pe26__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe26__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe26__lane31_strm1_data_mask   ;
  input                                           std__pe26__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe27__peId                ;
  input                                         sys__pe27__allSynchronized     ;
  output                                        pe27__sys__thisSynchronized    ;
  output                                        pe27__sys__ready               ;
  output                                        pe27__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe27__oob_cntl            ;
  input                                         std__pe27__oob_valid           ;
  output                                        pe27__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe27__oob_type            ;
  output                                          pe27__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane0_strm0_data_mask   ;
  input                                           std__pe27__lane0_strm0_data_valid  ;

  output                                          pe27__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane0_strm1_data_mask   ;
  input                                           std__pe27__lane0_strm1_data_valid  ;

  output                                          pe27__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane1_strm0_data_mask   ;
  input                                           std__pe27__lane1_strm0_data_valid  ;

  output                                          pe27__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane1_strm1_data_mask   ;
  input                                           std__pe27__lane1_strm1_data_valid  ;

  output                                          pe27__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane2_strm0_data_mask   ;
  input                                           std__pe27__lane2_strm0_data_valid  ;

  output                                          pe27__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane2_strm1_data_mask   ;
  input                                           std__pe27__lane2_strm1_data_valid  ;

  output                                          pe27__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane3_strm0_data_mask   ;
  input                                           std__pe27__lane3_strm0_data_valid  ;

  output                                          pe27__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane3_strm1_data_mask   ;
  input                                           std__pe27__lane3_strm1_data_valid  ;

  output                                          pe27__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane4_strm0_data_mask   ;
  input                                           std__pe27__lane4_strm0_data_valid  ;

  output                                          pe27__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane4_strm1_data_mask   ;
  input                                           std__pe27__lane4_strm1_data_valid  ;

  output                                          pe27__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane5_strm0_data_mask   ;
  input                                           std__pe27__lane5_strm0_data_valid  ;

  output                                          pe27__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane5_strm1_data_mask   ;
  input                                           std__pe27__lane5_strm1_data_valid  ;

  output                                          pe27__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane6_strm0_data_mask   ;
  input                                           std__pe27__lane6_strm0_data_valid  ;

  output                                          pe27__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane6_strm1_data_mask   ;
  input                                           std__pe27__lane6_strm1_data_valid  ;

  output                                          pe27__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane7_strm0_data_mask   ;
  input                                           std__pe27__lane7_strm0_data_valid  ;

  output                                          pe27__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane7_strm1_data_mask   ;
  input                                           std__pe27__lane7_strm1_data_valid  ;

  output                                          pe27__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane8_strm0_data_mask   ;
  input                                           std__pe27__lane8_strm0_data_valid  ;

  output                                          pe27__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane8_strm1_data_mask   ;
  input                                           std__pe27__lane8_strm1_data_valid  ;

  output                                          pe27__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane9_strm0_data_mask   ;
  input                                           std__pe27__lane9_strm0_data_valid  ;

  output                                          pe27__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane9_strm1_data_mask   ;
  input                                           std__pe27__lane9_strm1_data_valid  ;

  output                                          pe27__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane10_strm0_data_mask   ;
  input                                           std__pe27__lane10_strm0_data_valid  ;

  output                                          pe27__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane10_strm1_data_mask   ;
  input                                           std__pe27__lane10_strm1_data_valid  ;

  output                                          pe27__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane11_strm0_data_mask   ;
  input                                           std__pe27__lane11_strm0_data_valid  ;

  output                                          pe27__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane11_strm1_data_mask   ;
  input                                           std__pe27__lane11_strm1_data_valid  ;

  output                                          pe27__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane12_strm0_data_mask   ;
  input                                           std__pe27__lane12_strm0_data_valid  ;

  output                                          pe27__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane12_strm1_data_mask   ;
  input                                           std__pe27__lane12_strm1_data_valid  ;

  output                                          pe27__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane13_strm0_data_mask   ;
  input                                           std__pe27__lane13_strm0_data_valid  ;

  output                                          pe27__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane13_strm1_data_mask   ;
  input                                           std__pe27__lane13_strm1_data_valid  ;

  output                                          pe27__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane14_strm0_data_mask   ;
  input                                           std__pe27__lane14_strm0_data_valid  ;

  output                                          pe27__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane14_strm1_data_mask   ;
  input                                           std__pe27__lane14_strm1_data_valid  ;

  output                                          pe27__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane15_strm0_data_mask   ;
  input                                           std__pe27__lane15_strm0_data_valid  ;

  output                                          pe27__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane15_strm1_data_mask   ;
  input                                           std__pe27__lane15_strm1_data_valid  ;

  output                                          pe27__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane16_strm0_data_mask   ;
  input                                           std__pe27__lane16_strm0_data_valid  ;

  output                                          pe27__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane16_strm1_data_mask   ;
  input                                           std__pe27__lane16_strm1_data_valid  ;

  output                                          pe27__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane17_strm0_data_mask   ;
  input                                           std__pe27__lane17_strm0_data_valid  ;

  output                                          pe27__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane17_strm1_data_mask   ;
  input                                           std__pe27__lane17_strm1_data_valid  ;

  output                                          pe27__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane18_strm0_data_mask   ;
  input                                           std__pe27__lane18_strm0_data_valid  ;

  output                                          pe27__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane18_strm1_data_mask   ;
  input                                           std__pe27__lane18_strm1_data_valid  ;

  output                                          pe27__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane19_strm0_data_mask   ;
  input                                           std__pe27__lane19_strm0_data_valid  ;

  output                                          pe27__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane19_strm1_data_mask   ;
  input                                           std__pe27__lane19_strm1_data_valid  ;

  output                                          pe27__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane20_strm0_data_mask   ;
  input                                           std__pe27__lane20_strm0_data_valid  ;

  output                                          pe27__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane20_strm1_data_mask   ;
  input                                           std__pe27__lane20_strm1_data_valid  ;

  output                                          pe27__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane21_strm0_data_mask   ;
  input                                           std__pe27__lane21_strm0_data_valid  ;

  output                                          pe27__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane21_strm1_data_mask   ;
  input                                           std__pe27__lane21_strm1_data_valid  ;

  output                                          pe27__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane22_strm0_data_mask   ;
  input                                           std__pe27__lane22_strm0_data_valid  ;

  output                                          pe27__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane22_strm1_data_mask   ;
  input                                           std__pe27__lane22_strm1_data_valid  ;

  output                                          pe27__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane23_strm0_data_mask   ;
  input                                           std__pe27__lane23_strm0_data_valid  ;

  output                                          pe27__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane23_strm1_data_mask   ;
  input                                           std__pe27__lane23_strm1_data_valid  ;

  output                                          pe27__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane24_strm0_data_mask   ;
  input                                           std__pe27__lane24_strm0_data_valid  ;

  output                                          pe27__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane24_strm1_data_mask   ;
  input                                           std__pe27__lane24_strm1_data_valid  ;

  output                                          pe27__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane25_strm0_data_mask   ;
  input                                           std__pe27__lane25_strm0_data_valid  ;

  output                                          pe27__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane25_strm1_data_mask   ;
  input                                           std__pe27__lane25_strm1_data_valid  ;

  output                                          pe27__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane26_strm0_data_mask   ;
  input                                           std__pe27__lane26_strm0_data_valid  ;

  output                                          pe27__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane26_strm1_data_mask   ;
  input                                           std__pe27__lane26_strm1_data_valid  ;

  output                                          pe27__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane27_strm0_data_mask   ;
  input                                           std__pe27__lane27_strm0_data_valid  ;

  output                                          pe27__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane27_strm1_data_mask   ;
  input                                           std__pe27__lane27_strm1_data_valid  ;

  output                                          pe27__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane28_strm0_data_mask   ;
  input                                           std__pe27__lane28_strm0_data_valid  ;

  output                                          pe27__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane28_strm1_data_mask   ;
  input                                           std__pe27__lane28_strm1_data_valid  ;

  output                                          pe27__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane29_strm0_data_mask   ;
  input                                           std__pe27__lane29_strm0_data_valid  ;

  output                                          pe27__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane29_strm1_data_mask   ;
  input                                           std__pe27__lane29_strm1_data_valid  ;

  output                                          pe27__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane30_strm0_data_mask   ;
  input                                           std__pe27__lane30_strm0_data_valid  ;

  output                                          pe27__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane30_strm1_data_mask   ;
  input                                           std__pe27__lane30_strm1_data_valid  ;

  output                                          pe27__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane31_strm0_data_mask   ;
  input                                           std__pe27__lane31_strm0_data_valid  ;

  output                                          pe27__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe27__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe27__lane31_strm1_data_mask   ;
  input                                           std__pe27__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe28__peId                ;
  input                                         sys__pe28__allSynchronized     ;
  output                                        pe28__sys__thisSynchronized    ;
  output                                        pe28__sys__ready               ;
  output                                        pe28__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe28__oob_cntl            ;
  input                                         std__pe28__oob_valid           ;
  output                                        pe28__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe28__oob_type            ;
  output                                          pe28__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane0_strm0_data_mask   ;
  input                                           std__pe28__lane0_strm0_data_valid  ;

  output                                          pe28__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane0_strm1_data_mask   ;
  input                                           std__pe28__lane0_strm1_data_valid  ;

  output                                          pe28__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane1_strm0_data_mask   ;
  input                                           std__pe28__lane1_strm0_data_valid  ;

  output                                          pe28__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane1_strm1_data_mask   ;
  input                                           std__pe28__lane1_strm1_data_valid  ;

  output                                          pe28__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane2_strm0_data_mask   ;
  input                                           std__pe28__lane2_strm0_data_valid  ;

  output                                          pe28__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane2_strm1_data_mask   ;
  input                                           std__pe28__lane2_strm1_data_valid  ;

  output                                          pe28__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane3_strm0_data_mask   ;
  input                                           std__pe28__lane3_strm0_data_valid  ;

  output                                          pe28__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane3_strm1_data_mask   ;
  input                                           std__pe28__lane3_strm1_data_valid  ;

  output                                          pe28__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane4_strm0_data_mask   ;
  input                                           std__pe28__lane4_strm0_data_valid  ;

  output                                          pe28__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane4_strm1_data_mask   ;
  input                                           std__pe28__lane4_strm1_data_valid  ;

  output                                          pe28__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane5_strm0_data_mask   ;
  input                                           std__pe28__lane5_strm0_data_valid  ;

  output                                          pe28__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane5_strm1_data_mask   ;
  input                                           std__pe28__lane5_strm1_data_valid  ;

  output                                          pe28__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane6_strm0_data_mask   ;
  input                                           std__pe28__lane6_strm0_data_valid  ;

  output                                          pe28__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane6_strm1_data_mask   ;
  input                                           std__pe28__lane6_strm1_data_valid  ;

  output                                          pe28__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane7_strm0_data_mask   ;
  input                                           std__pe28__lane7_strm0_data_valid  ;

  output                                          pe28__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane7_strm1_data_mask   ;
  input                                           std__pe28__lane7_strm1_data_valid  ;

  output                                          pe28__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane8_strm0_data_mask   ;
  input                                           std__pe28__lane8_strm0_data_valid  ;

  output                                          pe28__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane8_strm1_data_mask   ;
  input                                           std__pe28__lane8_strm1_data_valid  ;

  output                                          pe28__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane9_strm0_data_mask   ;
  input                                           std__pe28__lane9_strm0_data_valid  ;

  output                                          pe28__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane9_strm1_data_mask   ;
  input                                           std__pe28__lane9_strm1_data_valid  ;

  output                                          pe28__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane10_strm0_data_mask   ;
  input                                           std__pe28__lane10_strm0_data_valid  ;

  output                                          pe28__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane10_strm1_data_mask   ;
  input                                           std__pe28__lane10_strm1_data_valid  ;

  output                                          pe28__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane11_strm0_data_mask   ;
  input                                           std__pe28__lane11_strm0_data_valid  ;

  output                                          pe28__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane11_strm1_data_mask   ;
  input                                           std__pe28__lane11_strm1_data_valid  ;

  output                                          pe28__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane12_strm0_data_mask   ;
  input                                           std__pe28__lane12_strm0_data_valid  ;

  output                                          pe28__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane12_strm1_data_mask   ;
  input                                           std__pe28__lane12_strm1_data_valid  ;

  output                                          pe28__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane13_strm0_data_mask   ;
  input                                           std__pe28__lane13_strm0_data_valid  ;

  output                                          pe28__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane13_strm1_data_mask   ;
  input                                           std__pe28__lane13_strm1_data_valid  ;

  output                                          pe28__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane14_strm0_data_mask   ;
  input                                           std__pe28__lane14_strm0_data_valid  ;

  output                                          pe28__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane14_strm1_data_mask   ;
  input                                           std__pe28__lane14_strm1_data_valid  ;

  output                                          pe28__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane15_strm0_data_mask   ;
  input                                           std__pe28__lane15_strm0_data_valid  ;

  output                                          pe28__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane15_strm1_data_mask   ;
  input                                           std__pe28__lane15_strm1_data_valid  ;

  output                                          pe28__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane16_strm0_data_mask   ;
  input                                           std__pe28__lane16_strm0_data_valid  ;

  output                                          pe28__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane16_strm1_data_mask   ;
  input                                           std__pe28__lane16_strm1_data_valid  ;

  output                                          pe28__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane17_strm0_data_mask   ;
  input                                           std__pe28__lane17_strm0_data_valid  ;

  output                                          pe28__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane17_strm1_data_mask   ;
  input                                           std__pe28__lane17_strm1_data_valid  ;

  output                                          pe28__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane18_strm0_data_mask   ;
  input                                           std__pe28__lane18_strm0_data_valid  ;

  output                                          pe28__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane18_strm1_data_mask   ;
  input                                           std__pe28__lane18_strm1_data_valid  ;

  output                                          pe28__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane19_strm0_data_mask   ;
  input                                           std__pe28__lane19_strm0_data_valid  ;

  output                                          pe28__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane19_strm1_data_mask   ;
  input                                           std__pe28__lane19_strm1_data_valid  ;

  output                                          pe28__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane20_strm0_data_mask   ;
  input                                           std__pe28__lane20_strm0_data_valid  ;

  output                                          pe28__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane20_strm1_data_mask   ;
  input                                           std__pe28__lane20_strm1_data_valid  ;

  output                                          pe28__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane21_strm0_data_mask   ;
  input                                           std__pe28__lane21_strm0_data_valid  ;

  output                                          pe28__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane21_strm1_data_mask   ;
  input                                           std__pe28__lane21_strm1_data_valid  ;

  output                                          pe28__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane22_strm0_data_mask   ;
  input                                           std__pe28__lane22_strm0_data_valid  ;

  output                                          pe28__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane22_strm1_data_mask   ;
  input                                           std__pe28__lane22_strm1_data_valid  ;

  output                                          pe28__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane23_strm0_data_mask   ;
  input                                           std__pe28__lane23_strm0_data_valid  ;

  output                                          pe28__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane23_strm1_data_mask   ;
  input                                           std__pe28__lane23_strm1_data_valid  ;

  output                                          pe28__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane24_strm0_data_mask   ;
  input                                           std__pe28__lane24_strm0_data_valid  ;

  output                                          pe28__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane24_strm1_data_mask   ;
  input                                           std__pe28__lane24_strm1_data_valid  ;

  output                                          pe28__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane25_strm0_data_mask   ;
  input                                           std__pe28__lane25_strm0_data_valid  ;

  output                                          pe28__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane25_strm1_data_mask   ;
  input                                           std__pe28__lane25_strm1_data_valid  ;

  output                                          pe28__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane26_strm0_data_mask   ;
  input                                           std__pe28__lane26_strm0_data_valid  ;

  output                                          pe28__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane26_strm1_data_mask   ;
  input                                           std__pe28__lane26_strm1_data_valid  ;

  output                                          pe28__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane27_strm0_data_mask   ;
  input                                           std__pe28__lane27_strm0_data_valid  ;

  output                                          pe28__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane27_strm1_data_mask   ;
  input                                           std__pe28__lane27_strm1_data_valid  ;

  output                                          pe28__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane28_strm0_data_mask   ;
  input                                           std__pe28__lane28_strm0_data_valid  ;

  output                                          pe28__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane28_strm1_data_mask   ;
  input                                           std__pe28__lane28_strm1_data_valid  ;

  output                                          pe28__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane29_strm0_data_mask   ;
  input                                           std__pe28__lane29_strm0_data_valid  ;

  output                                          pe28__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane29_strm1_data_mask   ;
  input                                           std__pe28__lane29_strm1_data_valid  ;

  output                                          pe28__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane30_strm0_data_mask   ;
  input                                           std__pe28__lane30_strm0_data_valid  ;

  output                                          pe28__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane30_strm1_data_mask   ;
  input                                           std__pe28__lane30_strm1_data_valid  ;

  output                                          pe28__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane31_strm0_data_mask   ;
  input                                           std__pe28__lane31_strm0_data_valid  ;

  output                                          pe28__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe28__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe28__lane31_strm1_data_mask   ;
  input                                           std__pe28__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe29__peId                ;
  input                                         sys__pe29__allSynchronized     ;
  output                                        pe29__sys__thisSynchronized    ;
  output                                        pe29__sys__ready               ;
  output                                        pe29__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe29__oob_cntl            ;
  input                                         std__pe29__oob_valid           ;
  output                                        pe29__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe29__oob_type            ;
  output                                          pe29__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane0_strm0_data_mask   ;
  input                                           std__pe29__lane0_strm0_data_valid  ;

  output                                          pe29__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane0_strm1_data_mask   ;
  input                                           std__pe29__lane0_strm1_data_valid  ;

  output                                          pe29__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane1_strm0_data_mask   ;
  input                                           std__pe29__lane1_strm0_data_valid  ;

  output                                          pe29__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane1_strm1_data_mask   ;
  input                                           std__pe29__lane1_strm1_data_valid  ;

  output                                          pe29__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane2_strm0_data_mask   ;
  input                                           std__pe29__lane2_strm0_data_valid  ;

  output                                          pe29__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane2_strm1_data_mask   ;
  input                                           std__pe29__lane2_strm1_data_valid  ;

  output                                          pe29__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane3_strm0_data_mask   ;
  input                                           std__pe29__lane3_strm0_data_valid  ;

  output                                          pe29__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane3_strm1_data_mask   ;
  input                                           std__pe29__lane3_strm1_data_valid  ;

  output                                          pe29__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane4_strm0_data_mask   ;
  input                                           std__pe29__lane4_strm0_data_valid  ;

  output                                          pe29__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane4_strm1_data_mask   ;
  input                                           std__pe29__lane4_strm1_data_valid  ;

  output                                          pe29__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane5_strm0_data_mask   ;
  input                                           std__pe29__lane5_strm0_data_valid  ;

  output                                          pe29__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane5_strm1_data_mask   ;
  input                                           std__pe29__lane5_strm1_data_valid  ;

  output                                          pe29__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane6_strm0_data_mask   ;
  input                                           std__pe29__lane6_strm0_data_valid  ;

  output                                          pe29__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane6_strm1_data_mask   ;
  input                                           std__pe29__lane6_strm1_data_valid  ;

  output                                          pe29__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane7_strm0_data_mask   ;
  input                                           std__pe29__lane7_strm0_data_valid  ;

  output                                          pe29__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane7_strm1_data_mask   ;
  input                                           std__pe29__lane7_strm1_data_valid  ;

  output                                          pe29__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane8_strm0_data_mask   ;
  input                                           std__pe29__lane8_strm0_data_valid  ;

  output                                          pe29__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane8_strm1_data_mask   ;
  input                                           std__pe29__lane8_strm1_data_valid  ;

  output                                          pe29__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane9_strm0_data_mask   ;
  input                                           std__pe29__lane9_strm0_data_valid  ;

  output                                          pe29__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane9_strm1_data_mask   ;
  input                                           std__pe29__lane9_strm1_data_valid  ;

  output                                          pe29__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane10_strm0_data_mask   ;
  input                                           std__pe29__lane10_strm0_data_valid  ;

  output                                          pe29__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane10_strm1_data_mask   ;
  input                                           std__pe29__lane10_strm1_data_valid  ;

  output                                          pe29__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane11_strm0_data_mask   ;
  input                                           std__pe29__lane11_strm0_data_valid  ;

  output                                          pe29__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane11_strm1_data_mask   ;
  input                                           std__pe29__lane11_strm1_data_valid  ;

  output                                          pe29__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane12_strm0_data_mask   ;
  input                                           std__pe29__lane12_strm0_data_valid  ;

  output                                          pe29__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane12_strm1_data_mask   ;
  input                                           std__pe29__lane12_strm1_data_valid  ;

  output                                          pe29__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane13_strm0_data_mask   ;
  input                                           std__pe29__lane13_strm0_data_valid  ;

  output                                          pe29__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane13_strm1_data_mask   ;
  input                                           std__pe29__lane13_strm1_data_valid  ;

  output                                          pe29__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane14_strm0_data_mask   ;
  input                                           std__pe29__lane14_strm0_data_valid  ;

  output                                          pe29__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane14_strm1_data_mask   ;
  input                                           std__pe29__lane14_strm1_data_valid  ;

  output                                          pe29__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane15_strm0_data_mask   ;
  input                                           std__pe29__lane15_strm0_data_valid  ;

  output                                          pe29__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane15_strm1_data_mask   ;
  input                                           std__pe29__lane15_strm1_data_valid  ;

  output                                          pe29__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane16_strm0_data_mask   ;
  input                                           std__pe29__lane16_strm0_data_valid  ;

  output                                          pe29__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane16_strm1_data_mask   ;
  input                                           std__pe29__lane16_strm1_data_valid  ;

  output                                          pe29__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane17_strm0_data_mask   ;
  input                                           std__pe29__lane17_strm0_data_valid  ;

  output                                          pe29__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane17_strm1_data_mask   ;
  input                                           std__pe29__lane17_strm1_data_valid  ;

  output                                          pe29__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane18_strm0_data_mask   ;
  input                                           std__pe29__lane18_strm0_data_valid  ;

  output                                          pe29__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane18_strm1_data_mask   ;
  input                                           std__pe29__lane18_strm1_data_valid  ;

  output                                          pe29__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane19_strm0_data_mask   ;
  input                                           std__pe29__lane19_strm0_data_valid  ;

  output                                          pe29__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane19_strm1_data_mask   ;
  input                                           std__pe29__lane19_strm1_data_valid  ;

  output                                          pe29__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane20_strm0_data_mask   ;
  input                                           std__pe29__lane20_strm0_data_valid  ;

  output                                          pe29__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane20_strm1_data_mask   ;
  input                                           std__pe29__lane20_strm1_data_valid  ;

  output                                          pe29__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane21_strm0_data_mask   ;
  input                                           std__pe29__lane21_strm0_data_valid  ;

  output                                          pe29__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane21_strm1_data_mask   ;
  input                                           std__pe29__lane21_strm1_data_valid  ;

  output                                          pe29__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane22_strm0_data_mask   ;
  input                                           std__pe29__lane22_strm0_data_valid  ;

  output                                          pe29__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane22_strm1_data_mask   ;
  input                                           std__pe29__lane22_strm1_data_valid  ;

  output                                          pe29__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane23_strm0_data_mask   ;
  input                                           std__pe29__lane23_strm0_data_valid  ;

  output                                          pe29__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane23_strm1_data_mask   ;
  input                                           std__pe29__lane23_strm1_data_valid  ;

  output                                          pe29__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane24_strm0_data_mask   ;
  input                                           std__pe29__lane24_strm0_data_valid  ;

  output                                          pe29__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane24_strm1_data_mask   ;
  input                                           std__pe29__lane24_strm1_data_valid  ;

  output                                          pe29__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane25_strm0_data_mask   ;
  input                                           std__pe29__lane25_strm0_data_valid  ;

  output                                          pe29__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane25_strm1_data_mask   ;
  input                                           std__pe29__lane25_strm1_data_valid  ;

  output                                          pe29__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane26_strm0_data_mask   ;
  input                                           std__pe29__lane26_strm0_data_valid  ;

  output                                          pe29__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane26_strm1_data_mask   ;
  input                                           std__pe29__lane26_strm1_data_valid  ;

  output                                          pe29__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane27_strm0_data_mask   ;
  input                                           std__pe29__lane27_strm0_data_valid  ;

  output                                          pe29__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane27_strm1_data_mask   ;
  input                                           std__pe29__lane27_strm1_data_valid  ;

  output                                          pe29__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane28_strm0_data_mask   ;
  input                                           std__pe29__lane28_strm0_data_valid  ;

  output                                          pe29__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane28_strm1_data_mask   ;
  input                                           std__pe29__lane28_strm1_data_valid  ;

  output                                          pe29__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane29_strm0_data_mask   ;
  input                                           std__pe29__lane29_strm0_data_valid  ;

  output                                          pe29__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane29_strm1_data_mask   ;
  input                                           std__pe29__lane29_strm1_data_valid  ;

  output                                          pe29__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane30_strm0_data_mask   ;
  input                                           std__pe29__lane30_strm0_data_valid  ;

  output                                          pe29__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane30_strm1_data_mask   ;
  input                                           std__pe29__lane30_strm1_data_valid  ;

  output                                          pe29__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane31_strm0_data_mask   ;
  input                                           std__pe29__lane31_strm0_data_valid  ;

  output                                          pe29__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe29__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe29__lane31_strm1_data_mask   ;
  input                                           std__pe29__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe30__peId                ;
  input                                         sys__pe30__allSynchronized     ;
  output                                        pe30__sys__thisSynchronized    ;
  output                                        pe30__sys__ready               ;
  output                                        pe30__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe30__oob_cntl            ;
  input                                         std__pe30__oob_valid           ;
  output                                        pe30__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe30__oob_type            ;
  output                                          pe30__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane0_strm0_data_mask   ;
  input                                           std__pe30__lane0_strm0_data_valid  ;

  output                                          pe30__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane0_strm1_data_mask   ;
  input                                           std__pe30__lane0_strm1_data_valid  ;

  output                                          pe30__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane1_strm0_data_mask   ;
  input                                           std__pe30__lane1_strm0_data_valid  ;

  output                                          pe30__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane1_strm1_data_mask   ;
  input                                           std__pe30__lane1_strm1_data_valid  ;

  output                                          pe30__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane2_strm0_data_mask   ;
  input                                           std__pe30__lane2_strm0_data_valid  ;

  output                                          pe30__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane2_strm1_data_mask   ;
  input                                           std__pe30__lane2_strm1_data_valid  ;

  output                                          pe30__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane3_strm0_data_mask   ;
  input                                           std__pe30__lane3_strm0_data_valid  ;

  output                                          pe30__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane3_strm1_data_mask   ;
  input                                           std__pe30__lane3_strm1_data_valid  ;

  output                                          pe30__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane4_strm0_data_mask   ;
  input                                           std__pe30__lane4_strm0_data_valid  ;

  output                                          pe30__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane4_strm1_data_mask   ;
  input                                           std__pe30__lane4_strm1_data_valid  ;

  output                                          pe30__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane5_strm0_data_mask   ;
  input                                           std__pe30__lane5_strm0_data_valid  ;

  output                                          pe30__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane5_strm1_data_mask   ;
  input                                           std__pe30__lane5_strm1_data_valid  ;

  output                                          pe30__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane6_strm0_data_mask   ;
  input                                           std__pe30__lane6_strm0_data_valid  ;

  output                                          pe30__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane6_strm1_data_mask   ;
  input                                           std__pe30__lane6_strm1_data_valid  ;

  output                                          pe30__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane7_strm0_data_mask   ;
  input                                           std__pe30__lane7_strm0_data_valid  ;

  output                                          pe30__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane7_strm1_data_mask   ;
  input                                           std__pe30__lane7_strm1_data_valid  ;

  output                                          pe30__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane8_strm0_data_mask   ;
  input                                           std__pe30__lane8_strm0_data_valid  ;

  output                                          pe30__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane8_strm1_data_mask   ;
  input                                           std__pe30__lane8_strm1_data_valid  ;

  output                                          pe30__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane9_strm0_data_mask   ;
  input                                           std__pe30__lane9_strm0_data_valid  ;

  output                                          pe30__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane9_strm1_data_mask   ;
  input                                           std__pe30__lane9_strm1_data_valid  ;

  output                                          pe30__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane10_strm0_data_mask   ;
  input                                           std__pe30__lane10_strm0_data_valid  ;

  output                                          pe30__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane10_strm1_data_mask   ;
  input                                           std__pe30__lane10_strm1_data_valid  ;

  output                                          pe30__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane11_strm0_data_mask   ;
  input                                           std__pe30__lane11_strm0_data_valid  ;

  output                                          pe30__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane11_strm1_data_mask   ;
  input                                           std__pe30__lane11_strm1_data_valid  ;

  output                                          pe30__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane12_strm0_data_mask   ;
  input                                           std__pe30__lane12_strm0_data_valid  ;

  output                                          pe30__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane12_strm1_data_mask   ;
  input                                           std__pe30__lane12_strm1_data_valid  ;

  output                                          pe30__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane13_strm0_data_mask   ;
  input                                           std__pe30__lane13_strm0_data_valid  ;

  output                                          pe30__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane13_strm1_data_mask   ;
  input                                           std__pe30__lane13_strm1_data_valid  ;

  output                                          pe30__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane14_strm0_data_mask   ;
  input                                           std__pe30__lane14_strm0_data_valid  ;

  output                                          pe30__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane14_strm1_data_mask   ;
  input                                           std__pe30__lane14_strm1_data_valid  ;

  output                                          pe30__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane15_strm0_data_mask   ;
  input                                           std__pe30__lane15_strm0_data_valid  ;

  output                                          pe30__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane15_strm1_data_mask   ;
  input                                           std__pe30__lane15_strm1_data_valid  ;

  output                                          pe30__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane16_strm0_data_mask   ;
  input                                           std__pe30__lane16_strm0_data_valid  ;

  output                                          pe30__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane16_strm1_data_mask   ;
  input                                           std__pe30__lane16_strm1_data_valid  ;

  output                                          pe30__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane17_strm0_data_mask   ;
  input                                           std__pe30__lane17_strm0_data_valid  ;

  output                                          pe30__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane17_strm1_data_mask   ;
  input                                           std__pe30__lane17_strm1_data_valid  ;

  output                                          pe30__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane18_strm0_data_mask   ;
  input                                           std__pe30__lane18_strm0_data_valid  ;

  output                                          pe30__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane18_strm1_data_mask   ;
  input                                           std__pe30__lane18_strm1_data_valid  ;

  output                                          pe30__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane19_strm0_data_mask   ;
  input                                           std__pe30__lane19_strm0_data_valid  ;

  output                                          pe30__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane19_strm1_data_mask   ;
  input                                           std__pe30__lane19_strm1_data_valid  ;

  output                                          pe30__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane20_strm0_data_mask   ;
  input                                           std__pe30__lane20_strm0_data_valid  ;

  output                                          pe30__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane20_strm1_data_mask   ;
  input                                           std__pe30__lane20_strm1_data_valid  ;

  output                                          pe30__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane21_strm0_data_mask   ;
  input                                           std__pe30__lane21_strm0_data_valid  ;

  output                                          pe30__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane21_strm1_data_mask   ;
  input                                           std__pe30__lane21_strm1_data_valid  ;

  output                                          pe30__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane22_strm0_data_mask   ;
  input                                           std__pe30__lane22_strm0_data_valid  ;

  output                                          pe30__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane22_strm1_data_mask   ;
  input                                           std__pe30__lane22_strm1_data_valid  ;

  output                                          pe30__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane23_strm0_data_mask   ;
  input                                           std__pe30__lane23_strm0_data_valid  ;

  output                                          pe30__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane23_strm1_data_mask   ;
  input                                           std__pe30__lane23_strm1_data_valid  ;

  output                                          pe30__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane24_strm0_data_mask   ;
  input                                           std__pe30__lane24_strm0_data_valid  ;

  output                                          pe30__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane24_strm1_data_mask   ;
  input                                           std__pe30__lane24_strm1_data_valid  ;

  output                                          pe30__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane25_strm0_data_mask   ;
  input                                           std__pe30__lane25_strm0_data_valid  ;

  output                                          pe30__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane25_strm1_data_mask   ;
  input                                           std__pe30__lane25_strm1_data_valid  ;

  output                                          pe30__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane26_strm0_data_mask   ;
  input                                           std__pe30__lane26_strm0_data_valid  ;

  output                                          pe30__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane26_strm1_data_mask   ;
  input                                           std__pe30__lane26_strm1_data_valid  ;

  output                                          pe30__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane27_strm0_data_mask   ;
  input                                           std__pe30__lane27_strm0_data_valid  ;

  output                                          pe30__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane27_strm1_data_mask   ;
  input                                           std__pe30__lane27_strm1_data_valid  ;

  output                                          pe30__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane28_strm0_data_mask   ;
  input                                           std__pe30__lane28_strm0_data_valid  ;

  output                                          pe30__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane28_strm1_data_mask   ;
  input                                           std__pe30__lane28_strm1_data_valid  ;

  output                                          pe30__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane29_strm0_data_mask   ;
  input                                           std__pe30__lane29_strm0_data_valid  ;

  output                                          pe30__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane29_strm1_data_mask   ;
  input                                           std__pe30__lane29_strm1_data_valid  ;

  output                                          pe30__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane30_strm0_data_mask   ;
  input                                           std__pe30__lane30_strm0_data_valid  ;

  output                                          pe30__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane30_strm1_data_mask   ;
  input                                           std__pe30__lane30_strm1_data_valid  ;

  output                                          pe30__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane31_strm0_data_mask   ;
  input                                           std__pe30__lane31_strm0_data_valid  ;

  output                                          pe30__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe30__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe30__lane31_strm1_data_mask   ;
  input                                           std__pe30__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe31__peId                ;
  input                                         sys__pe31__allSynchronized     ;
  output                                        pe31__sys__thisSynchronized    ;
  output                                        pe31__sys__ready               ;
  output                                        pe31__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe31__oob_cntl            ;
  input                                         std__pe31__oob_valid           ;
  output                                        pe31__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe31__oob_type            ;
  output                                          pe31__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane0_strm0_data_mask   ;
  input                                           std__pe31__lane0_strm0_data_valid  ;

  output                                          pe31__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane0_strm1_data_mask   ;
  input                                           std__pe31__lane0_strm1_data_valid  ;

  output                                          pe31__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane1_strm0_data_mask   ;
  input                                           std__pe31__lane1_strm0_data_valid  ;

  output                                          pe31__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane1_strm1_data_mask   ;
  input                                           std__pe31__lane1_strm1_data_valid  ;

  output                                          pe31__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane2_strm0_data_mask   ;
  input                                           std__pe31__lane2_strm0_data_valid  ;

  output                                          pe31__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane2_strm1_data_mask   ;
  input                                           std__pe31__lane2_strm1_data_valid  ;

  output                                          pe31__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane3_strm0_data_mask   ;
  input                                           std__pe31__lane3_strm0_data_valid  ;

  output                                          pe31__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane3_strm1_data_mask   ;
  input                                           std__pe31__lane3_strm1_data_valid  ;

  output                                          pe31__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane4_strm0_data_mask   ;
  input                                           std__pe31__lane4_strm0_data_valid  ;

  output                                          pe31__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane4_strm1_data_mask   ;
  input                                           std__pe31__lane4_strm1_data_valid  ;

  output                                          pe31__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane5_strm0_data_mask   ;
  input                                           std__pe31__lane5_strm0_data_valid  ;

  output                                          pe31__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane5_strm1_data_mask   ;
  input                                           std__pe31__lane5_strm1_data_valid  ;

  output                                          pe31__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane6_strm0_data_mask   ;
  input                                           std__pe31__lane6_strm0_data_valid  ;

  output                                          pe31__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane6_strm1_data_mask   ;
  input                                           std__pe31__lane6_strm1_data_valid  ;

  output                                          pe31__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane7_strm0_data_mask   ;
  input                                           std__pe31__lane7_strm0_data_valid  ;

  output                                          pe31__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane7_strm1_data_mask   ;
  input                                           std__pe31__lane7_strm1_data_valid  ;

  output                                          pe31__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane8_strm0_data_mask   ;
  input                                           std__pe31__lane8_strm0_data_valid  ;

  output                                          pe31__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane8_strm1_data_mask   ;
  input                                           std__pe31__lane8_strm1_data_valid  ;

  output                                          pe31__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane9_strm0_data_mask   ;
  input                                           std__pe31__lane9_strm0_data_valid  ;

  output                                          pe31__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane9_strm1_data_mask   ;
  input                                           std__pe31__lane9_strm1_data_valid  ;

  output                                          pe31__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane10_strm0_data_mask   ;
  input                                           std__pe31__lane10_strm0_data_valid  ;

  output                                          pe31__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane10_strm1_data_mask   ;
  input                                           std__pe31__lane10_strm1_data_valid  ;

  output                                          pe31__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane11_strm0_data_mask   ;
  input                                           std__pe31__lane11_strm0_data_valid  ;

  output                                          pe31__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane11_strm1_data_mask   ;
  input                                           std__pe31__lane11_strm1_data_valid  ;

  output                                          pe31__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane12_strm0_data_mask   ;
  input                                           std__pe31__lane12_strm0_data_valid  ;

  output                                          pe31__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane12_strm1_data_mask   ;
  input                                           std__pe31__lane12_strm1_data_valid  ;

  output                                          pe31__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane13_strm0_data_mask   ;
  input                                           std__pe31__lane13_strm0_data_valid  ;

  output                                          pe31__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane13_strm1_data_mask   ;
  input                                           std__pe31__lane13_strm1_data_valid  ;

  output                                          pe31__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane14_strm0_data_mask   ;
  input                                           std__pe31__lane14_strm0_data_valid  ;

  output                                          pe31__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane14_strm1_data_mask   ;
  input                                           std__pe31__lane14_strm1_data_valid  ;

  output                                          pe31__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane15_strm0_data_mask   ;
  input                                           std__pe31__lane15_strm0_data_valid  ;

  output                                          pe31__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane15_strm1_data_mask   ;
  input                                           std__pe31__lane15_strm1_data_valid  ;

  output                                          pe31__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane16_strm0_data_mask   ;
  input                                           std__pe31__lane16_strm0_data_valid  ;

  output                                          pe31__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane16_strm1_data_mask   ;
  input                                           std__pe31__lane16_strm1_data_valid  ;

  output                                          pe31__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane17_strm0_data_mask   ;
  input                                           std__pe31__lane17_strm0_data_valid  ;

  output                                          pe31__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane17_strm1_data_mask   ;
  input                                           std__pe31__lane17_strm1_data_valid  ;

  output                                          pe31__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane18_strm0_data_mask   ;
  input                                           std__pe31__lane18_strm0_data_valid  ;

  output                                          pe31__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane18_strm1_data_mask   ;
  input                                           std__pe31__lane18_strm1_data_valid  ;

  output                                          pe31__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane19_strm0_data_mask   ;
  input                                           std__pe31__lane19_strm0_data_valid  ;

  output                                          pe31__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane19_strm1_data_mask   ;
  input                                           std__pe31__lane19_strm1_data_valid  ;

  output                                          pe31__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane20_strm0_data_mask   ;
  input                                           std__pe31__lane20_strm0_data_valid  ;

  output                                          pe31__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane20_strm1_data_mask   ;
  input                                           std__pe31__lane20_strm1_data_valid  ;

  output                                          pe31__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane21_strm0_data_mask   ;
  input                                           std__pe31__lane21_strm0_data_valid  ;

  output                                          pe31__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane21_strm1_data_mask   ;
  input                                           std__pe31__lane21_strm1_data_valid  ;

  output                                          pe31__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane22_strm0_data_mask   ;
  input                                           std__pe31__lane22_strm0_data_valid  ;

  output                                          pe31__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane22_strm1_data_mask   ;
  input                                           std__pe31__lane22_strm1_data_valid  ;

  output                                          pe31__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane23_strm0_data_mask   ;
  input                                           std__pe31__lane23_strm0_data_valid  ;

  output                                          pe31__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane23_strm1_data_mask   ;
  input                                           std__pe31__lane23_strm1_data_valid  ;

  output                                          pe31__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane24_strm0_data_mask   ;
  input                                           std__pe31__lane24_strm0_data_valid  ;

  output                                          pe31__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane24_strm1_data_mask   ;
  input                                           std__pe31__lane24_strm1_data_valid  ;

  output                                          pe31__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane25_strm0_data_mask   ;
  input                                           std__pe31__lane25_strm0_data_valid  ;

  output                                          pe31__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane25_strm1_data_mask   ;
  input                                           std__pe31__lane25_strm1_data_valid  ;

  output                                          pe31__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane26_strm0_data_mask   ;
  input                                           std__pe31__lane26_strm0_data_valid  ;

  output                                          pe31__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane26_strm1_data_mask   ;
  input                                           std__pe31__lane26_strm1_data_valid  ;

  output                                          pe31__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane27_strm0_data_mask   ;
  input                                           std__pe31__lane27_strm0_data_valid  ;

  output                                          pe31__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane27_strm1_data_mask   ;
  input                                           std__pe31__lane27_strm1_data_valid  ;

  output                                          pe31__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane28_strm0_data_mask   ;
  input                                           std__pe31__lane28_strm0_data_valid  ;

  output                                          pe31__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane28_strm1_data_mask   ;
  input                                           std__pe31__lane28_strm1_data_valid  ;

  output                                          pe31__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane29_strm0_data_mask   ;
  input                                           std__pe31__lane29_strm0_data_valid  ;

  output                                          pe31__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane29_strm1_data_mask   ;
  input                                           std__pe31__lane29_strm1_data_valid  ;

  output                                          pe31__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane30_strm0_data_mask   ;
  input                                           std__pe31__lane30_strm0_data_valid  ;

  output                                          pe31__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane30_strm1_data_mask   ;
  input                                           std__pe31__lane30_strm1_data_valid  ;

  output                                          pe31__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane31_strm0_data_mask   ;
  input                                           std__pe31__lane31_strm0_data_valid  ;

  output                                          pe31__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe31__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe31__lane31_strm1_data_mask   ;
  input                                           std__pe31__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe32__peId                ;
  input                                         sys__pe32__allSynchronized     ;
  output                                        pe32__sys__thisSynchronized    ;
  output                                        pe32__sys__ready               ;
  output                                        pe32__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe32__oob_cntl            ;
  input                                         std__pe32__oob_valid           ;
  output                                        pe32__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe32__oob_type            ;
  output                                          pe32__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane0_strm0_data_mask   ;
  input                                           std__pe32__lane0_strm0_data_valid  ;

  output                                          pe32__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane0_strm1_data_mask   ;
  input                                           std__pe32__lane0_strm1_data_valid  ;

  output                                          pe32__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane1_strm0_data_mask   ;
  input                                           std__pe32__lane1_strm0_data_valid  ;

  output                                          pe32__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane1_strm1_data_mask   ;
  input                                           std__pe32__lane1_strm1_data_valid  ;

  output                                          pe32__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane2_strm0_data_mask   ;
  input                                           std__pe32__lane2_strm0_data_valid  ;

  output                                          pe32__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane2_strm1_data_mask   ;
  input                                           std__pe32__lane2_strm1_data_valid  ;

  output                                          pe32__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane3_strm0_data_mask   ;
  input                                           std__pe32__lane3_strm0_data_valid  ;

  output                                          pe32__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane3_strm1_data_mask   ;
  input                                           std__pe32__lane3_strm1_data_valid  ;

  output                                          pe32__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane4_strm0_data_mask   ;
  input                                           std__pe32__lane4_strm0_data_valid  ;

  output                                          pe32__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane4_strm1_data_mask   ;
  input                                           std__pe32__lane4_strm1_data_valid  ;

  output                                          pe32__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane5_strm0_data_mask   ;
  input                                           std__pe32__lane5_strm0_data_valid  ;

  output                                          pe32__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane5_strm1_data_mask   ;
  input                                           std__pe32__lane5_strm1_data_valid  ;

  output                                          pe32__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane6_strm0_data_mask   ;
  input                                           std__pe32__lane6_strm0_data_valid  ;

  output                                          pe32__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane6_strm1_data_mask   ;
  input                                           std__pe32__lane6_strm1_data_valid  ;

  output                                          pe32__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane7_strm0_data_mask   ;
  input                                           std__pe32__lane7_strm0_data_valid  ;

  output                                          pe32__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane7_strm1_data_mask   ;
  input                                           std__pe32__lane7_strm1_data_valid  ;

  output                                          pe32__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane8_strm0_data_mask   ;
  input                                           std__pe32__lane8_strm0_data_valid  ;

  output                                          pe32__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane8_strm1_data_mask   ;
  input                                           std__pe32__lane8_strm1_data_valid  ;

  output                                          pe32__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane9_strm0_data_mask   ;
  input                                           std__pe32__lane9_strm0_data_valid  ;

  output                                          pe32__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane9_strm1_data_mask   ;
  input                                           std__pe32__lane9_strm1_data_valid  ;

  output                                          pe32__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane10_strm0_data_mask   ;
  input                                           std__pe32__lane10_strm0_data_valid  ;

  output                                          pe32__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane10_strm1_data_mask   ;
  input                                           std__pe32__lane10_strm1_data_valid  ;

  output                                          pe32__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane11_strm0_data_mask   ;
  input                                           std__pe32__lane11_strm0_data_valid  ;

  output                                          pe32__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane11_strm1_data_mask   ;
  input                                           std__pe32__lane11_strm1_data_valid  ;

  output                                          pe32__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane12_strm0_data_mask   ;
  input                                           std__pe32__lane12_strm0_data_valid  ;

  output                                          pe32__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane12_strm1_data_mask   ;
  input                                           std__pe32__lane12_strm1_data_valid  ;

  output                                          pe32__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane13_strm0_data_mask   ;
  input                                           std__pe32__lane13_strm0_data_valid  ;

  output                                          pe32__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane13_strm1_data_mask   ;
  input                                           std__pe32__lane13_strm1_data_valid  ;

  output                                          pe32__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane14_strm0_data_mask   ;
  input                                           std__pe32__lane14_strm0_data_valid  ;

  output                                          pe32__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane14_strm1_data_mask   ;
  input                                           std__pe32__lane14_strm1_data_valid  ;

  output                                          pe32__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane15_strm0_data_mask   ;
  input                                           std__pe32__lane15_strm0_data_valid  ;

  output                                          pe32__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane15_strm1_data_mask   ;
  input                                           std__pe32__lane15_strm1_data_valid  ;

  output                                          pe32__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane16_strm0_data_mask   ;
  input                                           std__pe32__lane16_strm0_data_valid  ;

  output                                          pe32__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane16_strm1_data_mask   ;
  input                                           std__pe32__lane16_strm1_data_valid  ;

  output                                          pe32__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane17_strm0_data_mask   ;
  input                                           std__pe32__lane17_strm0_data_valid  ;

  output                                          pe32__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane17_strm1_data_mask   ;
  input                                           std__pe32__lane17_strm1_data_valid  ;

  output                                          pe32__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane18_strm0_data_mask   ;
  input                                           std__pe32__lane18_strm0_data_valid  ;

  output                                          pe32__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane18_strm1_data_mask   ;
  input                                           std__pe32__lane18_strm1_data_valid  ;

  output                                          pe32__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane19_strm0_data_mask   ;
  input                                           std__pe32__lane19_strm0_data_valid  ;

  output                                          pe32__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane19_strm1_data_mask   ;
  input                                           std__pe32__lane19_strm1_data_valid  ;

  output                                          pe32__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane20_strm0_data_mask   ;
  input                                           std__pe32__lane20_strm0_data_valid  ;

  output                                          pe32__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane20_strm1_data_mask   ;
  input                                           std__pe32__lane20_strm1_data_valid  ;

  output                                          pe32__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane21_strm0_data_mask   ;
  input                                           std__pe32__lane21_strm0_data_valid  ;

  output                                          pe32__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane21_strm1_data_mask   ;
  input                                           std__pe32__lane21_strm1_data_valid  ;

  output                                          pe32__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane22_strm0_data_mask   ;
  input                                           std__pe32__lane22_strm0_data_valid  ;

  output                                          pe32__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane22_strm1_data_mask   ;
  input                                           std__pe32__lane22_strm1_data_valid  ;

  output                                          pe32__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane23_strm0_data_mask   ;
  input                                           std__pe32__lane23_strm0_data_valid  ;

  output                                          pe32__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane23_strm1_data_mask   ;
  input                                           std__pe32__lane23_strm1_data_valid  ;

  output                                          pe32__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane24_strm0_data_mask   ;
  input                                           std__pe32__lane24_strm0_data_valid  ;

  output                                          pe32__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane24_strm1_data_mask   ;
  input                                           std__pe32__lane24_strm1_data_valid  ;

  output                                          pe32__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane25_strm0_data_mask   ;
  input                                           std__pe32__lane25_strm0_data_valid  ;

  output                                          pe32__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane25_strm1_data_mask   ;
  input                                           std__pe32__lane25_strm1_data_valid  ;

  output                                          pe32__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane26_strm0_data_mask   ;
  input                                           std__pe32__lane26_strm0_data_valid  ;

  output                                          pe32__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane26_strm1_data_mask   ;
  input                                           std__pe32__lane26_strm1_data_valid  ;

  output                                          pe32__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane27_strm0_data_mask   ;
  input                                           std__pe32__lane27_strm0_data_valid  ;

  output                                          pe32__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane27_strm1_data_mask   ;
  input                                           std__pe32__lane27_strm1_data_valid  ;

  output                                          pe32__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane28_strm0_data_mask   ;
  input                                           std__pe32__lane28_strm0_data_valid  ;

  output                                          pe32__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane28_strm1_data_mask   ;
  input                                           std__pe32__lane28_strm1_data_valid  ;

  output                                          pe32__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane29_strm0_data_mask   ;
  input                                           std__pe32__lane29_strm0_data_valid  ;

  output                                          pe32__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane29_strm1_data_mask   ;
  input                                           std__pe32__lane29_strm1_data_valid  ;

  output                                          pe32__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane30_strm0_data_mask   ;
  input                                           std__pe32__lane30_strm0_data_valid  ;

  output                                          pe32__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane30_strm1_data_mask   ;
  input                                           std__pe32__lane30_strm1_data_valid  ;

  output                                          pe32__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane31_strm0_data_mask   ;
  input                                           std__pe32__lane31_strm0_data_valid  ;

  output                                          pe32__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe32__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe32__lane31_strm1_data_mask   ;
  input                                           std__pe32__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe33__peId                ;
  input                                         sys__pe33__allSynchronized     ;
  output                                        pe33__sys__thisSynchronized    ;
  output                                        pe33__sys__ready               ;
  output                                        pe33__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe33__oob_cntl            ;
  input                                         std__pe33__oob_valid           ;
  output                                        pe33__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe33__oob_type            ;
  output                                          pe33__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane0_strm0_data_mask   ;
  input                                           std__pe33__lane0_strm0_data_valid  ;

  output                                          pe33__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane0_strm1_data_mask   ;
  input                                           std__pe33__lane0_strm1_data_valid  ;

  output                                          pe33__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane1_strm0_data_mask   ;
  input                                           std__pe33__lane1_strm0_data_valid  ;

  output                                          pe33__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane1_strm1_data_mask   ;
  input                                           std__pe33__lane1_strm1_data_valid  ;

  output                                          pe33__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane2_strm0_data_mask   ;
  input                                           std__pe33__lane2_strm0_data_valid  ;

  output                                          pe33__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane2_strm1_data_mask   ;
  input                                           std__pe33__lane2_strm1_data_valid  ;

  output                                          pe33__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane3_strm0_data_mask   ;
  input                                           std__pe33__lane3_strm0_data_valid  ;

  output                                          pe33__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane3_strm1_data_mask   ;
  input                                           std__pe33__lane3_strm1_data_valid  ;

  output                                          pe33__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane4_strm0_data_mask   ;
  input                                           std__pe33__lane4_strm0_data_valid  ;

  output                                          pe33__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane4_strm1_data_mask   ;
  input                                           std__pe33__lane4_strm1_data_valid  ;

  output                                          pe33__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane5_strm0_data_mask   ;
  input                                           std__pe33__lane5_strm0_data_valid  ;

  output                                          pe33__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane5_strm1_data_mask   ;
  input                                           std__pe33__lane5_strm1_data_valid  ;

  output                                          pe33__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane6_strm0_data_mask   ;
  input                                           std__pe33__lane6_strm0_data_valid  ;

  output                                          pe33__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane6_strm1_data_mask   ;
  input                                           std__pe33__lane6_strm1_data_valid  ;

  output                                          pe33__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane7_strm0_data_mask   ;
  input                                           std__pe33__lane7_strm0_data_valid  ;

  output                                          pe33__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane7_strm1_data_mask   ;
  input                                           std__pe33__lane7_strm1_data_valid  ;

  output                                          pe33__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane8_strm0_data_mask   ;
  input                                           std__pe33__lane8_strm0_data_valid  ;

  output                                          pe33__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane8_strm1_data_mask   ;
  input                                           std__pe33__lane8_strm1_data_valid  ;

  output                                          pe33__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane9_strm0_data_mask   ;
  input                                           std__pe33__lane9_strm0_data_valid  ;

  output                                          pe33__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane9_strm1_data_mask   ;
  input                                           std__pe33__lane9_strm1_data_valid  ;

  output                                          pe33__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane10_strm0_data_mask   ;
  input                                           std__pe33__lane10_strm0_data_valid  ;

  output                                          pe33__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane10_strm1_data_mask   ;
  input                                           std__pe33__lane10_strm1_data_valid  ;

  output                                          pe33__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane11_strm0_data_mask   ;
  input                                           std__pe33__lane11_strm0_data_valid  ;

  output                                          pe33__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane11_strm1_data_mask   ;
  input                                           std__pe33__lane11_strm1_data_valid  ;

  output                                          pe33__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane12_strm0_data_mask   ;
  input                                           std__pe33__lane12_strm0_data_valid  ;

  output                                          pe33__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane12_strm1_data_mask   ;
  input                                           std__pe33__lane12_strm1_data_valid  ;

  output                                          pe33__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane13_strm0_data_mask   ;
  input                                           std__pe33__lane13_strm0_data_valid  ;

  output                                          pe33__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane13_strm1_data_mask   ;
  input                                           std__pe33__lane13_strm1_data_valid  ;

  output                                          pe33__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane14_strm0_data_mask   ;
  input                                           std__pe33__lane14_strm0_data_valid  ;

  output                                          pe33__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane14_strm1_data_mask   ;
  input                                           std__pe33__lane14_strm1_data_valid  ;

  output                                          pe33__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane15_strm0_data_mask   ;
  input                                           std__pe33__lane15_strm0_data_valid  ;

  output                                          pe33__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane15_strm1_data_mask   ;
  input                                           std__pe33__lane15_strm1_data_valid  ;

  output                                          pe33__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane16_strm0_data_mask   ;
  input                                           std__pe33__lane16_strm0_data_valid  ;

  output                                          pe33__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane16_strm1_data_mask   ;
  input                                           std__pe33__lane16_strm1_data_valid  ;

  output                                          pe33__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane17_strm0_data_mask   ;
  input                                           std__pe33__lane17_strm0_data_valid  ;

  output                                          pe33__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane17_strm1_data_mask   ;
  input                                           std__pe33__lane17_strm1_data_valid  ;

  output                                          pe33__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane18_strm0_data_mask   ;
  input                                           std__pe33__lane18_strm0_data_valid  ;

  output                                          pe33__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane18_strm1_data_mask   ;
  input                                           std__pe33__lane18_strm1_data_valid  ;

  output                                          pe33__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane19_strm0_data_mask   ;
  input                                           std__pe33__lane19_strm0_data_valid  ;

  output                                          pe33__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane19_strm1_data_mask   ;
  input                                           std__pe33__lane19_strm1_data_valid  ;

  output                                          pe33__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane20_strm0_data_mask   ;
  input                                           std__pe33__lane20_strm0_data_valid  ;

  output                                          pe33__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane20_strm1_data_mask   ;
  input                                           std__pe33__lane20_strm1_data_valid  ;

  output                                          pe33__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane21_strm0_data_mask   ;
  input                                           std__pe33__lane21_strm0_data_valid  ;

  output                                          pe33__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane21_strm1_data_mask   ;
  input                                           std__pe33__lane21_strm1_data_valid  ;

  output                                          pe33__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane22_strm0_data_mask   ;
  input                                           std__pe33__lane22_strm0_data_valid  ;

  output                                          pe33__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane22_strm1_data_mask   ;
  input                                           std__pe33__lane22_strm1_data_valid  ;

  output                                          pe33__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane23_strm0_data_mask   ;
  input                                           std__pe33__lane23_strm0_data_valid  ;

  output                                          pe33__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane23_strm1_data_mask   ;
  input                                           std__pe33__lane23_strm1_data_valid  ;

  output                                          pe33__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane24_strm0_data_mask   ;
  input                                           std__pe33__lane24_strm0_data_valid  ;

  output                                          pe33__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane24_strm1_data_mask   ;
  input                                           std__pe33__lane24_strm1_data_valid  ;

  output                                          pe33__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane25_strm0_data_mask   ;
  input                                           std__pe33__lane25_strm0_data_valid  ;

  output                                          pe33__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane25_strm1_data_mask   ;
  input                                           std__pe33__lane25_strm1_data_valid  ;

  output                                          pe33__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane26_strm0_data_mask   ;
  input                                           std__pe33__lane26_strm0_data_valid  ;

  output                                          pe33__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane26_strm1_data_mask   ;
  input                                           std__pe33__lane26_strm1_data_valid  ;

  output                                          pe33__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane27_strm0_data_mask   ;
  input                                           std__pe33__lane27_strm0_data_valid  ;

  output                                          pe33__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane27_strm1_data_mask   ;
  input                                           std__pe33__lane27_strm1_data_valid  ;

  output                                          pe33__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane28_strm0_data_mask   ;
  input                                           std__pe33__lane28_strm0_data_valid  ;

  output                                          pe33__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane28_strm1_data_mask   ;
  input                                           std__pe33__lane28_strm1_data_valid  ;

  output                                          pe33__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane29_strm0_data_mask   ;
  input                                           std__pe33__lane29_strm0_data_valid  ;

  output                                          pe33__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane29_strm1_data_mask   ;
  input                                           std__pe33__lane29_strm1_data_valid  ;

  output                                          pe33__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane30_strm0_data_mask   ;
  input                                           std__pe33__lane30_strm0_data_valid  ;

  output                                          pe33__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane30_strm1_data_mask   ;
  input                                           std__pe33__lane30_strm1_data_valid  ;

  output                                          pe33__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane31_strm0_data_mask   ;
  input                                           std__pe33__lane31_strm0_data_valid  ;

  output                                          pe33__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe33__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe33__lane31_strm1_data_mask   ;
  input                                           std__pe33__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe34__peId                ;
  input                                         sys__pe34__allSynchronized     ;
  output                                        pe34__sys__thisSynchronized    ;
  output                                        pe34__sys__ready               ;
  output                                        pe34__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe34__oob_cntl            ;
  input                                         std__pe34__oob_valid           ;
  output                                        pe34__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe34__oob_type            ;
  output                                          pe34__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane0_strm0_data_mask   ;
  input                                           std__pe34__lane0_strm0_data_valid  ;

  output                                          pe34__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane0_strm1_data_mask   ;
  input                                           std__pe34__lane0_strm1_data_valid  ;

  output                                          pe34__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane1_strm0_data_mask   ;
  input                                           std__pe34__lane1_strm0_data_valid  ;

  output                                          pe34__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane1_strm1_data_mask   ;
  input                                           std__pe34__lane1_strm1_data_valid  ;

  output                                          pe34__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane2_strm0_data_mask   ;
  input                                           std__pe34__lane2_strm0_data_valid  ;

  output                                          pe34__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane2_strm1_data_mask   ;
  input                                           std__pe34__lane2_strm1_data_valid  ;

  output                                          pe34__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane3_strm0_data_mask   ;
  input                                           std__pe34__lane3_strm0_data_valid  ;

  output                                          pe34__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane3_strm1_data_mask   ;
  input                                           std__pe34__lane3_strm1_data_valid  ;

  output                                          pe34__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane4_strm0_data_mask   ;
  input                                           std__pe34__lane4_strm0_data_valid  ;

  output                                          pe34__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane4_strm1_data_mask   ;
  input                                           std__pe34__lane4_strm1_data_valid  ;

  output                                          pe34__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane5_strm0_data_mask   ;
  input                                           std__pe34__lane5_strm0_data_valid  ;

  output                                          pe34__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane5_strm1_data_mask   ;
  input                                           std__pe34__lane5_strm1_data_valid  ;

  output                                          pe34__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane6_strm0_data_mask   ;
  input                                           std__pe34__lane6_strm0_data_valid  ;

  output                                          pe34__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane6_strm1_data_mask   ;
  input                                           std__pe34__lane6_strm1_data_valid  ;

  output                                          pe34__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane7_strm0_data_mask   ;
  input                                           std__pe34__lane7_strm0_data_valid  ;

  output                                          pe34__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane7_strm1_data_mask   ;
  input                                           std__pe34__lane7_strm1_data_valid  ;

  output                                          pe34__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane8_strm0_data_mask   ;
  input                                           std__pe34__lane8_strm0_data_valid  ;

  output                                          pe34__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane8_strm1_data_mask   ;
  input                                           std__pe34__lane8_strm1_data_valid  ;

  output                                          pe34__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane9_strm0_data_mask   ;
  input                                           std__pe34__lane9_strm0_data_valid  ;

  output                                          pe34__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane9_strm1_data_mask   ;
  input                                           std__pe34__lane9_strm1_data_valid  ;

  output                                          pe34__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane10_strm0_data_mask   ;
  input                                           std__pe34__lane10_strm0_data_valid  ;

  output                                          pe34__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane10_strm1_data_mask   ;
  input                                           std__pe34__lane10_strm1_data_valid  ;

  output                                          pe34__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane11_strm0_data_mask   ;
  input                                           std__pe34__lane11_strm0_data_valid  ;

  output                                          pe34__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane11_strm1_data_mask   ;
  input                                           std__pe34__lane11_strm1_data_valid  ;

  output                                          pe34__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane12_strm0_data_mask   ;
  input                                           std__pe34__lane12_strm0_data_valid  ;

  output                                          pe34__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane12_strm1_data_mask   ;
  input                                           std__pe34__lane12_strm1_data_valid  ;

  output                                          pe34__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane13_strm0_data_mask   ;
  input                                           std__pe34__lane13_strm0_data_valid  ;

  output                                          pe34__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane13_strm1_data_mask   ;
  input                                           std__pe34__lane13_strm1_data_valid  ;

  output                                          pe34__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane14_strm0_data_mask   ;
  input                                           std__pe34__lane14_strm0_data_valid  ;

  output                                          pe34__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane14_strm1_data_mask   ;
  input                                           std__pe34__lane14_strm1_data_valid  ;

  output                                          pe34__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane15_strm0_data_mask   ;
  input                                           std__pe34__lane15_strm0_data_valid  ;

  output                                          pe34__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane15_strm1_data_mask   ;
  input                                           std__pe34__lane15_strm1_data_valid  ;

  output                                          pe34__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane16_strm0_data_mask   ;
  input                                           std__pe34__lane16_strm0_data_valid  ;

  output                                          pe34__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane16_strm1_data_mask   ;
  input                                           std__pe34__lane16_strm1_data_valid  ;

  output                                          pe34__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane17_strm0_data_mask   ;
  input                                           std__pe34__lane17_strm0_data_valid  ;

  output                                          pe34__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane17_strm1_data_mask   ;
  input                                           std__pe34__lane17_strm1_data_valid  ;

  output                                          pe34__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane18_strm0_data_mask   ;
  input                                           std__pe34__lane18_strm0_data_valid  ;

  output                                          pe34__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane18_strm1_data_mask   ;
  input                                           std__pe34__lane18_strm1_data_valid  ;

  output                                          pe34__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane19_strm0_data_mask   ;
  input                                           std__pe34__lane19_strm0_data_valid  ;

  output                                          pe34__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane19_strm1_data_mask   ;
  input                                           std__pe34__lane19_strm1_data_valid  ;

  output                                          pe34__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane20_strm0_data_mask   ;
  input                                           std__pe34__lane20_strm0_data_valid  ;

  output                                          pe34__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane20_strm1_data_mask   ;
  input                                           std__pe34__lane20_strm1_data_valid  ;

  output                                          pe34__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane21_strm0_data_mask   ;
  input                                           std__pe34__lane21_strm0_data_valid  ;

  output                                          pe34__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane21_strm1_data_mask   ;
  input                                           std__pe34__lane21_strm1_data_valid  ;

  output                                          pe34__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane22_strm0_data_mask   ;
  input                                           std__pe34__lane22_strm0_data_valid  ;

  output                                          pe34__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane22_strm1_data_mask   ;
  input                                           std__pe34__lane22_strm1_data_valid  ;

  output                                          pe34__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane23_strm0_data_mask   ;
  input                                           std__pe34__lane23_strm0_data_valid  ;

  output                                          pe34__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane23_strm1_data_mask   ;
  input                                           std__pe34__lane23_strm1_data_valid  ;

  output                                          pe34__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane24_strm0_data_mask   ;
  input                                           std__pe34__lane24_strm0_data_valid  ;

  output                                          pe34__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane24_strm1_data_mask   ;
  input                                           std__pe34__lane24_strm1_data_valid  ;

  output                                          pe34__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane25_strm0_data_mask   ;
  input                                           std__pe34__lane25_strm0_data_valid  ;

  output                                          pe34__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane25_strm1_data_mask   ;
  input                                           std__pe34__lane25_strm1_data_valid  ;

  output                                          pe34__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane26_strm0_data_mask   ;
  input                                           std__pe34__lane26_strm0_data_valid  ;

  output                                          pe34__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane26_strm1_data_mask   ;
  input                                           std__pe34__lane26_strm1_data_valid  ;

  output                                          pe34__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane27_strm0_data_mask   ;
  input                                           std__pe34__lane27_strm0_data_valid  ;

  output                                          pe34__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane27_strm1_data_mask   ;
  input                                           std__pe34__lane27_strm1_data_valid  ;

  output                                          pe34__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane28_strm0_data_mask   ;
  input                                           std__pe34__lane28_strm0_data_valid  ;

  output                                          pe34__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane28_strm1_data_mask   ;
  input                                           std__pe34__lane28_strm1_data_valid  ;

  output                                          pe34__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane29_strm0_data_mask   ;
  input                                           std__pe34__lane29_strm0_data_valid  ;

  output                                          pe34__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane29_strm1_data_mask   ;
  input                                           std__pe34__lane29_strm1_data_valid  ;

  output                                          pe34__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane30_strm0_data_mask   ;
  input                                           std__pe34__lane30_strm0_data_valid  ;

  output                                          pe34__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane30_strm1_data_mask   ;
  input                                           std__pe34__lane30_strm1_data_valid  ;

  output                                          pe34__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane31_strm0_data_mask   ;
  input                                           std__pe34__lane31_strm0_data_valid  ;

  output                                          pe34__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe34__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe34__lane31_strm1_data_mask   ;
  input                                           std__pe34__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe35__peId                ;
  input                                         sys__pe35__allSynchronized     ;
  output                                        pe35__sys__thisSynchronized    ;
  output                                        pe35__sys__ready               ;
  output                                        pe35__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe35__oob_cntl            ;
  input                                         std__pe35__oob_valid           ;
  output                                        pe35__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe35__oob_type            ;
  output                                          pe35__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane0_strm0_data_mask   ;
  input                                           std__pe35__lane0_strm0_data_valid  ;

  output                                          pe35__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane0_strm1_data_mask   ;
  input                                           std__pe35__lane0_strm1_data_valid  ;

  output                                          pe35__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane1_strm0_data_mask   ;
  input                                           std__pe35__lane1_strm0_data_valid  ;

  output                                          pe35__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane1_strm1_data_mask   ;
  input                                           std__pe35__lane1_strm1_data_valid  ;

  output                                          pe35__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane2_strm0_data_mask   ;
  input                                           std__pe35__lane2_strm0_data_valid  ;

  output                                          pe35__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane2_strm1_data_mask   ;
  input                                           std__pe35__lane2_strm1_data_valid  ;

  output                                          pe35__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane3_strm0_data_mask   ;
  input                                           std__pe35__lane3_strm0_data_valid  ;

  output                                          pe35__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane3_strm1_data_mask   ;
  input                                           std__pe35__lane3_strm1_data_valid  ;

  output                                          pe35__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane4_strm0_data_mask   ;
  input                                           std__pe35__lane4_strm0_data_valid  ;

  output                                          pe35__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane4_strm1_data_mask   ;
  input                                           std__pe35__lane4_strm1_data_valid  ;

  output                                          pe35__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane5_strm0_data_mask   ;
  input                                           std__pe35__lane5_strm0_data_valid  ;

  output                                          pe35__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane5_strm1_data_mask   ;
  input                                           std__pe35__lane5_strm1_data_valid  ;

  output                                          pe35__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane6_strm0_data_mask   ;
  input                                           std__pe35__lane6_strm0_data_valid  ;

  output                                          pe35__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane6_strm1_data_mask   ;
  input                                           std__pe35__lane6_strm1_data_valid  ;

  output                                          pe35__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane7_strm0_data_mask   ;
  input                                           std__pe35__lane7_strm0_data_valid  ;

  output                                          pe35__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane7_strm1_data_mask   ;
  input                                           std__pe35__lane7_strm1_data_valid  ;

  output                                          pe35__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane8_strm0_data_mask   ;
  input                                           std__pe35__lane8_strm0_data_valid  ;

  output                                          pe35__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane8_strm1_data_mask   ;
  input                                           std__pe35__lane8_strm1_data_valid  ;

  output                                          pe35__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane9_strm0_data_mask   ;
  input                                           std__pe35__lane9_strm0_data_valid  ;

  output                                          pe35__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane9_strm1_data_mask   ;
  input                                           std__pe35__lane9_strm1_data_valid  ;

  output                                          pe35__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane10_strm0_data_mask   ;
  input                                           std__pe35__lane10_strm0_data_valid  ;

  output                                          pe35__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane10_strm1_data_mask   ;
  input                                           std__pe35__lane10_strm1_data_valid  ;

  output                                          pe35__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane11_strm0_data_mask   ;
  input                                           std__pe35__lane11_strm0_data_valid  ;

  output                                          pe35__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane11_strm1_data_mask   ;
  input                                           std__pe35__lane11_strm1_data_valid  ;

  output                                          pe35__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane12_strm0_data_mask   ;
  input                                           std__pe35__lane12_strm0_data_valid  ;

  output                                          pe35__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane12_strm1_data_mask   ;
  input                                           std__pe35__lane12_strm1_data_valid  ;

  output                                          pe35__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane13_strm0_data_mask   ;
  input                                           std__pe35__lane13_strm0_data_valid  ;

  output                                          pe35__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane13_strm1_data_mask   ;
  input                                           std__pe35__lane13_strm1_data_valid  ;

  output                                          pe35__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane14_strm0_data_mask   ;
  input                                           std__pe35__lane14_strm0_data_valid  ;

  output                                          pe35__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane14_strm1_data_mask   ;
  input                                           std__pe35__lane14_strm1_data_valid  ;

  output                                          pe35__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane15_strm0_data_mask   ;
  input                                           std__pe35__lane15_strm0_data_valid  ;

  output                                          pe35__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane15_strm1_data_mask   ;
  input                                           std__pe35__lane15_strm1_data_valid  ;

  output                                          pe35__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane16_strm0_data_mask   ;
  input                                           std__pe35__lane16_strm0_data_valid  ;

  output                                          pe35__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane16_strm1_data_mask   ;
  input                                           std__pe35__lane16_strm1_data_valid  ;

  output                                          pe35__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane17_strm0_data_mask   ;
  input                                           std__pe35__lane17_strm0_data_valid  ;

  output                                          pe35__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane17_strm1_data_mask   ;
  input                                           std__pe35__lane17_strm1_data_valid  ;

  output                                          pe35__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane18_strm0_data_mask   ;
  input                                           std__pe35__lane18_strm0_data_valid  ;

  output                                          pe35__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane18_strm1_data_mask   ;
  input                                           std__pe35__lane18_strm1_data_valid  ;

  output                                          pe35__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane19_strm0_data_mask   ;
  input                                           std__pe35__lane19_strm0_data_valid  ;

  output                                          pe35__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane19_strm1_data_mask   ;
  input                                           std__pe35__lane19_strm1_data_valid  ;

  output                                          pe35__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane20_strm0_data_mask   ;
  input                                           std__pe35__lane20_strm0_data_valid  ;

  output                                          pe35__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane20_strm1_data_mask   ;
  input                                           std__pe35__lane20_strm1_data_valid  ;

  output                                          pe35__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane21_strm0_data_mask   ;
  input                                           std__pe35__lane21_strm0_data_valid  ;

  output                                          pe35__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane21_strm1_data_mask   ;
  input                                           std__pe35__lane21_strm1_data_valid  ;

  output                                          pe35__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane22_strm0_data_mask   ;
  input                                           std__pe35__lane22_strm0_data_valid  ;

  output                                          pe35__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane22_strm1_data_mask   ;
  input                                           std__pe35__lane22_strm1_data_valid  ;

  output                                          pe35__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane23_strm0_data_mask   ;
  input                                           std__pe35__lane23_strm0_data_valid  ;

  output                                          pe35__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane23_strm1_data_mask   ;
  input                                           std__pe35__lane23_strm1_data_valid  ;

  output                                          pe35__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane24_strm0_data_mask   ;
  input                                           std__pe35__lane24_strm0_data_valid  ;

  output                                          pe35__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane24_strm1_data_mask   ;
  input                                           std__pe35__lane24_strm1_data_valid  ;

  output                                          pe35__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane25_strm0_data_mask   ;
  input                                           std__pe35__lane25_strm0_data_valid  ;

  output                                          pe35__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane25_strm1_data_mask   ;
  input                                           std__pe35__lane25_strm1_data_valid  ;

  output                                          pe35__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane26_strm0_data_mask   ;
  input                                           std__pe35__lane26_strm0_data_valid  ;

  output                                          pe35__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane26_strm1_data_mask   ;
  input                                           std__pe35__lane26_strm1_data_valid  ;

  output                                          pe35__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane27_strm0_data_mask   ;
  input                                           std__pe35__lane27_strm0_data_valid  ;

  output                                          pe35__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane27_strm1_data_mask   ;
  input                                           std__pe35__lane27_strm1_data_valid  ;

  output                                          pe35__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane28_strm0_data_mask   ;
  input                                           std__pe35__lane28_strm0_data_valid  ;

  output                                          pe35__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane28_strm1_data_mask   ;
  input                                           std__pe35__lane28_strm1_data_valid  ;

  output                                          pe35__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane29_strm0_data_mask   ;
  input                                           std__pe35__lane29_strm0_data_valid  ;

  output                                          pe35__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane29_strm1_data_mask   ;
  input                                           std__pe35__lane29_strm1_data_valid  ;

  output                                          pe35__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane30_strm0_data_mask   ;
  input                                           std__pe35__lane30_strm0_data_valid  ;

  output                                          pe35__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane30_strm1_data_mask   ;
  input                                           std__pe35__lane30_strm1_data_valid  ;

  output                                          pe35__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane31_strm0_data_mask   ;
  input                                           std__pe35__lane31_strm0_data_valid  ;

  output                                          pe35__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe35__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe35__lane31_strm1_data_mask   ;
  input                                           std__pe35__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe36__peId                ;
  input                                         sys__pe36__allSynchronized     ;
  output                                        pe36__sys__thisSynchronized    ;
  output                                        pe36__sys__ready               ;
  output                                        pe36__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe36__oob_cntl            ;
  input                                         std__pe36__oob_valid           ;
  output                                        pe36__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe36__oob_type            ;
  output                                          pe36__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane0_strm0_data_mask   ;
  input                                           std__pe36__lane0_strm0_data_valid  ;

  output                                          pe36__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane0_strm1_data_mask   ;
  input                                           std__pe36__lane0_strm1_data_valid  ;

  output                                          pe36__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane1_strm0_data_mask   ;
  input                                           std__pe36__lane1_strm0_data_valid  ;

  output                                          pe36__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane1_strm1_data_mask   ;
  input                                           std__pe36__lane1_strm1_data_valid  ;

  output                                          pe36__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane2_strm0_data_mask   ;
  input                                           std__pe36__lane2_strm0_data_valid  ;

  output                                          pe36__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane2_strm1_data_mask   ;
  input                                           std__pe36__lane2_strm1_data_valid  ;

  output                                          pe36__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane3_strm0_data_mask   ;
  input                                           std__pe36__lane3_strm0_data_valid  ;

  output                                          pe36__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane3_strm1_data_mask   ;
  input                                           std__pe36__lane3_strm1_data_valid  ;

  output                                          pe36__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane4_strm0_data_mask   ;
  input                                           std__pe36__lane4_strm0_data_valid  ;

  output                                          pe36__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane4_strm1_data_mask   ;
  input                                           std__pe36__lane4_strm1_data_valid  ;

  output                                          pe36__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane5_strm0_data_mask   ;
  input                                           std__pe36__lane5_strm0_data_valid  ;

  output                                          pe36__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane5_strm1_data_mask   ;
  input                                           std__pe36__lane5_strm1_data_valid  ;

  output                                          pe36__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane6_strm0_data_mask   ;
  input                                           std__pe36__lane6_strm0_data_valid  ;

  output                                          pe36__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane6_strm1_data_mask   ;
  input                                           std__pe36__lane6_strm1_data_valid  ;

  output                                          pe36__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane7_strm0_data_mask   ;
  input                                           std__pe36__lane7_strm0_data_valid  ;

  output                                          pe36__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane7_strm1_data_mask   ;
  input                                           std__pe36__lane7_strm1_data_valid  ;

  output                                          pe36__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane8_strm0_data_mask   ;
  input                                           std__pe36__lane8_strm0_data_valid  ;

  output                                          pe36__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane8_strm1_data_mask   ;
  input                                           std__pe36__lane8_strm1_data_valid  ;

  output                                          pe36__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane9_strm0_data_mask   ;
  input                                           std__pe36__lane9_strm0_data_valid  ;

  output                                          pe36__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane9_strm1_data_mask   ;
  input                                           std__pe36__lane9_strm1_data_valid  ;

  output                                          pe36__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane10_strm0_data_mask   ;
  input                                           std__pe36__lane10_strm0_data_valid  ;

  output                                          pe36__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane10_strm1_data_mask   ;
  input                                           std__pe36__lane10_strm1_data_valid  ;

  output                                          pe36__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane11_strm0_data_mask   ;
  input                                           std__pe36__lane11_strm0_data_valid  ;

  output                                          pe36__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane11_strm1_data_mask   ;
  input                                           std__pe36__lane11_strm1_data_valid  ;

  output                                          pe36__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane12_strm0_data_mask   ;
  input                                           std__pe36__lane12_strm0_data_valid  ;

  output                                          pe36__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane12_strm1_data_mask   ;
  input                                           std__pe36__lane12_strm1_data_valid  ;

  output                                          pe36__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane13_strm0_data_mask   ;
  input                                           std__pe36__lane13_strm0_data_valid  ;

  output                                          pe36__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane13_strm1_data_mask   ;
  input                                           std__pe36__lane13_strm1_data_valid  ;

  output                                          pe36__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane14_strm0_data_mask   ;
  input                                           std__pe36__lane14_strm0_data_valid  ;

  output                                          pe36__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane14_strm1_data_mask   ;
  input                                           std__pe36__lane14_strm1_data_valid  ;

  output                                          pe36__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane15_strm0_data_mask   ;
  input                                           std__pe36__lane15_strm0_data_valid  ;

  output                                          pe36__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane15_strm1_data_mask   ;
  input                                           std__pe36__lane15_strm1_data_valid  ;

  output                                          pe36__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane16_strm0_data_mask   ;
  input                                           std__pe36__lane16_strm0_data_valid  ;

  output                                          pe36__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane16_strm1_data_mask   ;
  input                                           std__pe36__lane16_strm1_data_valid  ;

  output                                          pe36__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane17_strm0_data_mask   ;
  input                                           std__pe36__lane17_strm0_data_valid  ;

  output                                          pe36__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane17_strm1_data_mask   ;
  input                                           std__pe36__lane17_strm1_data_valid  ;

  output                                          pe36__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane18_strm0_data_mask   ;
  input                                           std__pe36__lane18_strm0_data_valid  ;

  output                                          pe36__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane18_strm1_data_mask   ;
  input                                           std__pe36__lane18_strm1_data_valid  ;

  output                                          pe36__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane19_strm0_data_mask   ;
  input                                           std__pe36__lane19_strm0_data_valid  ;

  output                                          pe36__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane19_strm1_data_mask   ;
  input                                           std__pe36__lane19_strm1_data_valid  ;

  output                                          pe36__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane20_strm0_data_mask   ;
  input                                           std__pe36__lane20_strm0_data_valid  ;

  output                                          pe36__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane20_strm1_data_mask   ;
  input                                           std__pe36__lane20_strm1_data_valid  ;

  output                                          pe36__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane21_strm0_data_mask   ;
  input                                           std__pe36__lane21_strm0_data_valid  ;

  output                                          pe36__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane21_strm1_data_mask   ;
  input                                           std__pe36__lane21_strm1_data_valid  ;

  output                                          pe36__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane22_strm0_data_mask   ;
  input                                           std__pe36__lane22_strm0_data_valid  ;

  output                                          pe36__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane22_strm1_data_mask   ;
  input                                           std__pe36__lane22_strm1_data_valid  ;

  output                                          pe36__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane23_strm0_data_mask   ;
  input                                           std__pe36__lane23_strm0_data_valid  ;

  output                                          pe36__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane23_strm1_data_mask   ;
  input                                           std__pe36__lane23_strm1_data_valid  ;

  output                                          pe36__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane24_strm0_data_mask   ;
  input                                           std__pe36__lane24_strm0_data_valid  ;

  output                                          pe36__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane24_strm1_data_mask   ;
  input                                           std__pe36__lane24_strm1_data_valid  ;

  output                                          pe36__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane25_strm0_data_mask   ;
  input                                           std__pe36__lane25_strm0_data_valid  ;

  output                                          pe36__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane25_strm1_data_mask   ;
  input                                           std__pe36__lane25_strm1_data_valid  ;

  output                                          pe36__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane26_strm0_data_mask   ;
  input                                           std__pe36__lane26_strm0_data_valid  ;

  output                                          pe36__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane26_strm1_data_mask   ;
  input                                           std__pe36__lane26_strm1_data_valid  ;

  output                                          pe36__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane27_strm0_data_mask   ;
  input                                           std__pe36__lane27_strm0_data_valid  ;

  output                                          pe36__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane27_strm1_data_mask   ;
  input                                           std__pe36__lane27_strm1_data_valid  ;

  output                                          pe36__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane28_strm0_data_mask   ;
  input                                           std__pe36__lane28_strm0_data_valid  ;

  output                                          pe36__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane28_strm1_data_mask   ;
  input                                           std__pe36__lane28_strm1_data_valid  ;

  output                                          pe36__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane29_strm0_data_mask   ;
  input                                           std__pe36__lane29_strm0_data_valid  ;

  output                                          pe36__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane29_strm1_data_mask   ;
  input                                           std__pe36__lane29_strm1_data_valid  ;

  output                                          pe36__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane30_strm0_data_mask   ;
  input                                           std__pe36__lane30_strm0_data_valid  ;

  output                                          pe36__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane30_strm1_data_mask   ;
  input                                           std__pe36__lane30_strm1_data_valid  ;

  output                                          pe36__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane31_strm0_data_mask   ;
  input                                           std__pe36__lane31_strm0_data_valid  ;

  output                                          pe36__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe36__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe36__lane31_strm1_data_mask   ;
  input                                           std__pe36__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe37__peId                ;
  input                                         sys__pe37__allSynchronized     ;
  output                                        pe37__sys__thisSynchronized    ;
  output                                        pe37__sys__ready               ;
  output                                        pe37__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe37__oob_cntl            ;
  input                                         std__pe37__oob_valid           ;
  output                                        pe37__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe37__oob_type            ;
  output                                          pe37__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane0_strm0_data_mask   ;
  input                                           std__pe37__lane0_strm0_data_valid  ;

  output                                          pe37__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane0_strm1_data_mask   ;
  input                                           std__pe37__lane0_strm1_data_valid  ;

  output                                          pe37__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane1_strm0_data_mask   ;
  input                                           std__pe37__lane1_strm0_data_valid  ;

  output                                          pe37__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane1_strm1_data_mask   ;
  input                                           std__pe37__lane1_strm1_data_valid  ;

  output                                          pe37__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane2_strm0_data_mask   ;
  input                                           std__pe37__lane2_strm0_data_valid  ;

  output                                          pe37__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane2_strm1_data_mask   ;
  input                                           std__pe37__lane2_strm1_data_valid  ;

  output                                          pe37__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane3_strm0_data_mask   ;
  input                                           std__pe37__lane3_strm0_data_valid  ;

  output                                          pe37__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane3_strm1_data_mask   ;
  input                                           std__pe37__lane3_strm1_data_valid  ;

  output                                          pe37__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane4_strm0_data_mask   ;
  input                                           std__pe37__lane4_strm0_data_valid  ;

  output                                          pe37__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane4_strm1_data_mask   ;
  input                                           std__pe37__lane4_strm1_data_valid  ;

  output                                          pe37__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane5_strm0_data_mask   ;
  input                                           std__pe37__lane5_strm0_data_valid  ;

  output                                          pe37__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane5_strm1_data_mask   ;
  input                                           std__pe37__lane5_strm1_data_valid  ;

  output                                          pe37__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane6_strm0_data_mask   ;
  input                                           std__pe37__lane6_strm0_data_valid  ;

  output                                          pe37__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane6_strm1_data_mask   ;
  input                                           std__pe37__lane6_strm1_data_valid  ;

  output                                          pe37__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane7_strm0_data_mask   ;
  input                                           std__pe37__lane7_strm0_data_valid  ;

  output                                          pe37__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane7_strm1_data_mask   ;
  input                                           std__pe37__lane7_strm1_data_valid  ;

  output                                          pe37__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane8_strm0_data_mask   ;
  input                                           std__pe37__lane8_strm0_data_valid  ;

  output                                          pe37__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane8_strm1_data_mask   ;
  input                                           std__pe37__lane8_strm1_data_valid  ;

  output                                          pe37__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane9_strm0_data_mask   ;
  input                                           std__pe37__lane9_strm0_data_valid  ;

  output                                          pe37__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane9_strm1_data_mask   ;
  input                                           std__pe37__lane9_strm1_data_valid  ;

  output                                          pe37__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane10_strm0_data_mask   ;
  input                                           std__pe37__lane10_strm0_data_valid  ;

  output                                          pe37__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane10_strm1_data_mask   ;
  input                                           std__pe37__lane10_strm1_data_valid  ;

  output                                          pe37__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane11_strm0_data_mask   ;
  input                                           std__pe37__lane11_strm0_data_valid  ;

  output                                          pe37__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane11_strm1_data_mask   ;
  input                                           std__pe37__lane11_strm1_data_valid  ;

  output                                          pe37__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane12_strm0_data_mask   ;
  input                                           std__pe37__lane12_strm0_data_valid  ;

  output                                          pe37__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane12_strm1_data_mask   ;
  input                                           std__pe37__lane12_strm1_data_valid  ;

  output                                          pe37__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane13_strm0_data_mask   ;
  input                                           std__pe37__lane13_strm0_data_valid  ;

  output                                          pe37__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane13_strm1_data_mask   ;
  input                                           std__pe37__lane13_strm1_data_valid  ;

  output                                          pe37__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane14_strm0_data_mask   ;
  input                                           std__pe37__lane14_strm0_data_valid  ;

  output                                          pe37__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane14_strm1_data_mask   ;
  input                                           std__pe37__lane14_strm1_data_valid  ;

  output                                          pe37__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane15_strm0_data_mask   ;
  input                                           std__pe37__lane15_strm0_data_valid  ;

  output                                          pe37__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane15_strm1_data_mask   ;
  input                                           std__pe37__lane15_strm1_data_valid  ;

  output                                          pe37__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane16_strm0_data_mask   ;
  input                                           std__pe37__lane16_strm0_data_valid  ;

  output                                          pe37__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane16_strm1_data_mask   ;
  input                                           std__pe37__lane16_strm1_data_valid  ;

  output                                          pe37__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane17_strm0_data_mask   ;
  input                                           std__pe37__lane17_strm0_data_valid  ;

  output                                          pe37__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane17_strm1_data_mask   ;
  input                                           std__pe37__lane17_strm1_data_valid  ;

  output                                          pe37__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane18_strm0_data_mask   ;
  input                                           std__pe37__lane18_strm0_data_valid  ;

  output                                          pe37__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane18_strm1_data_mask   ;
  input                                           std__pe37__lane18_strm1_data_valid  ;

  output                                          pe37__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane19_strm0_data_mask   ;
  input                                           std__pe37__lane19_strm0_data_valid  ;

  output                                          pe37__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane19_strm1_data_mask   ;
  input                                           std__pe37__lane19_strm1_data_valid  ;

  output                                          pe37__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane20_strm0_data_mask   ;
  input                                           std__pe37__lane20_strm0_data_valid  ;

  output                                          pe37__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane20_strm1_data_mask   ;
  input                                           std__pe37__lane20_strm1_data_valid  ;

  output                                          pe37__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane21_strm0_data_mask   ;
  input                                           std__pe37__lane21_strm0_data_valid  ;

  output                                          pe37__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane21_strm1_data_mask   ;
  input                                           std__pe37__lane21_strm1_data_valid  ;

  output                                          pe37__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane22_strm0_data_mask   ;
  input                                           std__pe37__lane22_strm0_data_valid  ;

  output                                          pe37__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane22_strm1_data_mask   ;
  input                                           std__pe37__lane22_strm1_data_valid  ;

  output                                          pe37__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane23_strm0_data_mask   ;
  input                                           std__pe37__lane23_strm0_data_valid  ;

  output                                          pe37__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane23_strm1_data_mask   ;
  input                                           std__pe37__lane23_strm1_data_valid  ;

  output                                          pe37__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane24_strm0_data_mask   ;
  input                                           std__pe37__lane24_strm0_data_valid  ;

  output                                          pe37__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane24_strm1_data_mask   ;
  input                                           std__pe37__lane24_strm1_data_valid  ;

  output                                          pe37__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane25_strm0_data_mask   ;
  input                                           std__pe37__lane25_strm0_data_valid  ;

  output                                          pe37__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane25_strm1_data_mask   ;
  input                                           std__pe37__lane25_strm1_data_valid  ;

  output                                          pe37__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane26_strm0_data_mask   ;
  input                                           std__pe37__lane26_strm0_data_valid  ;

  output                                          pe37__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane26_strm1_data_mask   ;
  input                                           std__pe37__lane26_strm1_data_valid  ;

  output                                          pe37__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane27_strm0_data_mask   ;
  input                                           std__pe37__lane27_strm0_data_valid  ;

  output                                          pe37__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane27_strm1_data_mask   ;
  input                                           std__pe37__lane27_strm1_data_valid  ;

  output                                          pe37__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane28_strm0_data_mask   ;
  input                                           std__pe37__lane28_strm0_data_valid  ;

  output                                          pe37__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane28_strm1_data_mask   ;
  input                                           std__pe37__lane28_strm1_data_valid  ;

  output                                          pe37__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane29_strm0_data_mask   ;
  input                                           std__pe37__lane29_strm0_data_valid  ;

  output                                          pe37__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane29_strm1_data_mask   ;
  input                                           std__pe37__lane29_strm1_data_valid  ;

  output                                          pe37__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane30_strm0_data_mask   ;
  input                                           std__pe37__lane30_strm0_data_valid  ;

  output                                          pe37__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane30_strm1_data_mask   ;
  input                                           std__pe37__lane30_strm1_data_valid  ;

  output                                          pe37__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane31_strm0_data_mask   ;
  input                                           std__pe37__lane31_strm0_data_valid  ;

  output                                          pe37__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe37__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe37__lane31_strm1_data_mask   ;
  input                                           std__pe37__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe38__peId                ;
  input                                         sys__pe38__allSynchronized     ;
  output                                        pe38__sys__thisSynchronized    ;
  output                                        pe38__sys__ready               ;
  output                                        pe38__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe38__oob_cntl            ;
  input                                         std__pe38__oob_valid           ;
  output                                        pe38__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe38__oob_type            ;
  output                                          pe38__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane0_strm0_data_mask   ;
  input                                           std__pe38__lane0_strm0_data_valid  ;

  output                                          pe38__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane0_strm1_data_mask   ;
  input                                           std__pe38__lane0_strm1_data_valid  ;

  output                                          pe38__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane1_strm0_data_mask   ;
  input                                           std__pe38__lane1_strm0_data_valid  ;

  output                                          pe38__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane1_strm1_data_mask   ;
  input                                           std__pe38__lane1_strm1_data_valid  ;

  output                                          pe38__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane2_strm0_data_mask   ;
  input                                           std__pe38__lane2_strm0_data_valid  ;

  output                                          pe38__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane2_strm1_data_mask   ;
  input                                           std__pe38__lane2_strm1_data_valid  ;

  output                                          pe38__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane3_strm0_data_mask   ;
  input                                           std__pe38__lane3_strm0_data_valid  ;

  output                                          pe38__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane3_strm1_data_mask   ;
  input                                           std__pe38__lane3_strm1_data_valid  ;

  output                                          pe38__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane4_strm0_data_mask   ;
  input                                           std__pe38__lane4_strm0_data_valid  ;

  output                                          pe38__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane4_strm1_data_mask   ;
  input                                           std__pe38__lane4_strm1_data_valid  ;

  output                                          pe38__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane5_strm0_data_mask   ;
  input                                           std__pe38__lane5_strm0_data_valid  ;

  output                                          pe38__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane5_strm1_data_mask   ;
  input                                           std__pe38__lane5_strm1_data_valid  ;

  output                                          pe38__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane6_strm0_data_mask   ;
  input                                           std__pe38__lane6_strm0_data_valid  ;

  output                                          pe38__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane6_strm1_data_mask   ;
  input                                           std__pe38__lane6_strm1_data_valid  ;

  output                                          pe38__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane7_strm0_data_mask   ;
  input                                           std__pe38__lane7_strm0_data_valid  ;

  output                                          pe38__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane7_strm1_data_mask   ;
  input                                           std__pe38__lane7_strm1_data_valid  ;

  output                                          pe38__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane8_strm0_data_mask   ;
  input                                           std__pe38__lane8_strm0_data_valid  ;

  output                                          pe38__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane8_strm1_data_mask   ;
  input                                           std__pe38__lane8_strm1_data_valid  ;

  output                                          pe38__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane9_strm0_data_mask   ;
  input                                           std__pe38__lane9_strm0_data_valid  ;

  output                                          pe38__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane9_strm1_data_mask   ;
  input                                           std__pe38__lane9_strm1_data_valid  ;

  output                                          pe38__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane10_strm0_data_mask   ;
  input                                           std__pe38__lane10_strm0_data_valid  ;

  output                                          pe38__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane10_strm1_data_mask   ;
  input                                           std__pe38__lane10_strm1_data_valid  ;

  output                                          pe38__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane11_strm0_data_mask   ;
  input                                           std__pe38__lane11_strm0_data_valid  ;

  output                                          pe38__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane11_strm1_data_mask   ;
  input                                           std__pe38__lane11_strm1_data_valid  ;

  output                                          pe38__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane12_strm0_data_mask   ;
  input                                           std__pe38__lane12_strm0_data_valid  ;

  output                                          pe38__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane12_strm1_data_mask   ;
  input                                           std__pe38__lane12_strm1_data_valid  ;

  output                                          pe38__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane13_strm0_data_mask   ;
  input                                           std__pe38__lane13_strm0_data_valid  ;

  output                                          pe38__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane13_strm1_data_mask   ;
  input                                           std__pe38__lane13_strm1_data_valid  ;

  output                                          pe38__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane14_strm0_data_mask   ;
  input                                           std__pe38__lane14_strm0_data_valid  ;

  output                                          pe38__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane14_strm1_data_mask   ;
  input                                           std__pe38__lane14_strm1_data_valid  ;

  output                                          pe38__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane15_strm0_data_mask   ;
  input                                           std__pe38__lane15_strm0_data_valid  ;

  output                                          pe38__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane15_strm1_data_mask   ;
  input                                           std__pe38__lane15_strm1_data_valid  ;

  output                                          pe38__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane16_strm0_data_mask   ;
  input                                           std__pe38__lane16_strm0_data_valid  ;

  output                                          pe38__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane16_strm1_data_mask   ;
  input                                           std__pe38__lane16_strm1_data_valid  ;

  output                                          pe38__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane17_strm0_data_mask   ;
  input                                           std__pe38__lane17_strm0_data_valid  ;

  output                                          pe38__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane17_strm1_data_mask   ;
  input                                           std__pe38__lane17_strm1_data_valid  ;

  output                                          pe38__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane18_strm0_data_mask   ;
  input                                           std__pe38__lane18_strm0_data_valid  ;

  output                                          pe38__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane18_strm1_data_mask   ;
  input                                           std__pe38__lane18_strm1_data_valid  ;

  output                                          pe38__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane19_strm0_data_mask   ;
  input                                           std__pe38__lane19_strm0_data_valid  ;

  output                                          pe38__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane19_strm1_data_mask   ;
  input                                           std__pe38__lane19_strm1_data_valid  ;

  output                                          pe38__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane20_strm0_data_mask   ;
  input                                           std__pe38__lane20_strm0_data_valid  ;

  output                                          pe38__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane20_strm1_data_mask   ;
  input                                           std__pe38__lane20_strm1_data_valid  ;

  output                                          pe38__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane21_strm0_data_mask   ;
  input                                           std__pe38__lane21_strm0_data_valid  ;

  output                                          pe38__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane21_strm1_data_mask   ;
  input                                           std__pe38__lane21_strm1_data_valid  ;

  output                                          pe38__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane22_strm0_data_mask   ;
  input                                           std__pe38__lane22_strm0_data_valid  ;

  output                                          pe38__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane22_strm1_data_mask   ;
  input                                           std__pe38__lane22_strm1_data_valid  ;

  output                                          pe38__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane23_strm0_data_mask   ;
  input                                           std__pe38__lane23_strm0_data_valid  ;

  output                                          pe38__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane23_strm1_data_mask   ;
  input                                           std__pe38__lane23_strm1_data_valid  ;

  output                                          pe38__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane24_strm0_data_mask   ;
  input                                           std__pe38__lane24_strm0_data_valid  ;

  output                                          pe38__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane24_strm1_data_mask   ;
  input                                           std__pe38__lane24_strm1_data_valid  ;

  output                                          pe38__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane25_strm0_data_mask   ;
  input                                           std__pe38__lane25_strm0_data_valid  ;

  output                                          pe38__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane25_strm1_data_mask   ;
  input                                           std__pe38__lane25_strm1_data_valid  ;

  output                                          pe38__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane26_strm0_data_mask   ;
  input                                           std__pe38__lane26_strm0_data_valid  ;

  output                                          pe38__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane26_strm1_data_mask   ;
  input                                           std__pe38__lane26_strm1_data_valid  ;

  output                                          pe38__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane27_strm0_data_mask   ;
  input                                           std__pe38__lane27_strm0_data_valid  ;

  output                                          pe38__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane27_strm1_data_mask   ;
  input                                           std__pe38__lane27_strm1_data_valid  ;

  output                                          pe38__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane28_strm0_data_mask   ;
  input                                           std__pe38__lane28_strm0_data_valid  ;

  output                                          pe38__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane28_strm1_data_mask   ;
  input                                           std__pe38__lane28_strm1_data_valid  ;

  output                                          pe38__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane29_strm0_data_mask   ;
  input                                           std__pe38__lane29_strm0_data_valid  ;

  output                                          pe38__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane29_strm1_data_mask   ;
  input                                           std__pe38__lane29_strm1_data_valid  ;

  output                                          pe38__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane30_strm0_data_mask   ;
  input                                           std__pe38__lane30_strm0_data_valid  ;

  output                                          pe38__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane30_strm1_data_mask   ;
  input                                           std__pe38__lane30_strm1_data_valid  ;

  output                                          pe38__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane31_strm0_data_mask   ;
  input                                           std__pe38__lane31_strm0_data_valid  ;

  output                                          pe38__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe38__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe38__lane31_strm1_data_mask   ;
  input                                           std__pe38__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe39__peId                ;
  input                                         sys__pe39__allSynchronized     ;
  output                                        pe39__sys__thisSynchronized    ;
  output                                        pe39__sys__ready               ;
  output                                        pe39__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe39__oob_cntl            ;
  input                                         std__pe39__oob_valid           ;
  output                                        pe39__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe39__oob_type            ;
  output                                          pe39__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane0_strm0_data_mask   ;
  input                                           std__pe39__lane0_strm0_data_valid  ;

  output                                          pe39__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane0_strm1_data_mask   ;
  input                                           std__pe39__lane0_strm1_data_valid  ;

  output                                          pe39__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane1_strm0_data_mask   ;
  input                                           std__pe39__lane1_strm0_data_valid  ;

  output                                          pe39__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane1_strm1_data_mask   ;
  input                                           std__pe39__lane1_strm1_data_valid  ;

  output                                          pe39__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane2_strm0_data_mask   ;
  input                                           std__pe39__lane2_strm0_data_valid  ;

  output                                          pe39__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane2_strm1_data_mask   ;
  input                                           std__pe39__lane2_strm1_data_valid  ;

  output                                          pe39__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane3_strm0_data_mask   ;
  input                                           std__pe39__lane3_strm0_data_valid  ;

  output                                          pe39__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane3_strm1_data_mask   ;
  input                                           std__pe39__lane3_strm1_data_valid  ;

  output                                          pe39__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane4_strm0_data_mask   ;
  input                                           std__pe39__lane4_strm0_data_valid  ;

  output                                          pe39__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane4_strm1_data_mask   ;
  input                                           std__pe39__lane4_strm1_data_valid  ;

  output                                          pe39__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane5_strm0_data_mask   ;
  input                                           std__pe39__lane5_strm0_data_valid  ;

  output                                          pe39__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane5_strm1_data_mask   ;
  input                                           std__pe39__lane5_strm1_data_valid  ;

  output                                          pe39__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane6_strm0_data_mask   ;
  input                                           std__pe39__lane6_strm0_data_valid  ;

  output                                          pe39__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane6_strm1_data_mask   ;
  input                                           std__pe39__lane6_strm1_data_valid  ;

  output                                          pe39__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane7_strm0_data_mask   ;
  input                                           std__pe39__lane7_strm0_data_valid  ;

  output                                          pe39__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane7_strm1_data_mask   ;
  input                                           std__pe39__lane7_strm1_data_valid  ;

  output                                          pe39__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane8_strm0_data_mask   ;
  input                                           std__pe39__lane8_strm0_data_valid  ;

  output                                          pe39__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane8_strm1_data_mask   ;
  input                                           std__pe39__lane8_strm1_data_valid  ;

  output                                          pe39__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane9_strm0_data_mask   ;
  input                                           std__pe39__lane9_strm0_data_valid  ;

  output                                          pe39__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane9_strm1_data_mask   ;
  input                                           std__pe39__lane9_strm1_data_valid  ;

  output                                          pe39__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane10_strm0_data_mask   ;
  input                                           std__pe39__lane10_strm0_data_valid  ;

  output                                          pe39__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane10_strm1_data_mask   ;
  input                                           std__pe39__lane10_strm1_data_valid  ;

  output                                          pe39__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane11_strm0_data_mask   ;
  input                                           std__pe39__lane11_strm0_data_valid  ;

  output                                          pe39__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane11_strm1_data_mask   ;
  input                                           std__pe39__lane11_strm1_data_valid  ;

  output                                          pe39__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane12_strm0_data_mask   ;
  input                                           std__pe39__lane12_strm0_data_valid  ;

  output                                          pe39__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane12_strm1_data_mask   ;
  input                                           std__pe39__lane12_strm1_data_valid  ;

  output                                          pe39__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane13_strm0_data_mask   ;
  input                                           std__pe39__lane13_strm0_data_valid  ;

  output                                          pe39__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane13_strm1_data_mask   ;
  input                                           std__pe39__lane13_strm1_data_valid  ;

  output                                          pe39__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane14_strm0_data_mask   ;
  input                                           std__pe39__lane14_strm0_data_valid  ;

  output                                          pe39__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane14_strm1_data_mask   ;
  input                                           std__pe39__lane14_strm1_data_valid  ;

  output                                          pe39__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane15_strm0_data_mask   ;
  input                                           std__pe39__lane15_strm0_data_valid  ;

  output                                          pe39__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane15_strm1_data_mask   ;
  input                                           std__pe39__lane15_strm1_data_valid  ;

  output                                          pe39__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane16_strm0_data_mask   ;
  input                                           std__pe39__lane16_strm0_data_valid  ;

  output                                          pe39__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane16_strm1_data_mask   ;
  input                                           std__pe39__lane16_strm1_data_valid  ;

  output                                          pe39__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane17_strm0_data_mask   ;
  input                                           std__pe39__lane17_strm0_data_valid  ;

  output                                          pe39__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane17_strm1_data_mask   ;
  input                                           std__pe39__lane17_strm1_data_valid  ;

  output                                          pe39__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane18_strm0_data_mask   ;
  input                                           std__pe39__lane18_strm0_data_valid  ;

  output                                          pe39__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane18_strm1_data_mask   ;
  input                                           std__pe39__lane18_strm1_data_valid  ;

  output                                          pe39__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane19_strm0_data_mask   ;
  input                                           std__pe39__lane19_strm0_data_valid  ;

  output                                          pe39__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane19_strm1_data_mask   ;
  input                                           std__pe39__lane19_strm1_data_valid  ;

  output                                          pe39__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane20_strm0_data_mask   ;
  input                                           std__pe39__lane20_strm0_data_valid  ;

  output                                          pe39__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane20_strm1_data_mask   ;
  input                                           std__pe39__lane20_strm1_data_valid  ;

  output                                          pe39__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane21_strm0_data_mask   ;
  input                                           std__pe39__lane21_strm0_data_valid  ;

  output                                          pe39__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane21_strm1_data_mask   ;
  input                                           std__pe39__lane21_strm1_data_valid  ;

  output                                          pe39__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane22_strm0_data_mask   ;
  input                                           std__pe39__lane22_strm0_data_valid  ;

  output                                          pe39__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane22_strm1_data_mask   ;
  input                                           std__pe39__lane22_strm1_data_valid  ;

  output                                          pe39__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane23_strm0_data_mask   ;
  input                                           std__pe39__lane23_strm0_data_valid  ;

  output                                          pe39__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane23_strm1_data_mask   ;
  input                                           std__pe39__lane23_strm1_data_valid  ;

  output                                          pe39__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane24_strm0_data_mask   ;
  input                                           std__pe39__lane24_strm0_data_valid  ;

  output                                          pe39__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane24_strm1_data_mask   ;
  input                                           std__pe39__lane24_strm1_data_valid  ;

  output                                          pe39__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane25_strm0_data_mask   ;
  input                                           std__pe39__lane25_strm0_data_valid  ;

  output                                          pe39__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane25_strm1_data_mask   ;
  input                                           std__pe39__lane25_strm1_data_valid  ;

  output                                          pe39__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane26_strm0_data_mask   ;
  input                                           std__pe39__lane26_strm0_data_valid  ;

  output                                          pe39__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane26_strm1_data_mask   ;
  input                                           std__pe39__lane26_strm1_data_valid  ;

  output                                          pe39__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane27_strm0_data_mask   ;
  input                                           std__pe39__lane27_strm0_data_valid  ;

  output                                          pe39__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane27_strm1_data_mask   ;
  input                                           std__pe39__lane27_strm1_data_valid  ;

  output                                          pe39__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane28_strm0_data_mask   ;
  input                                           std__pe39__lane28_strm0_data_valid  ;

  output                                          pe39__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane28_strm1_data_mask   ;
  input                                           std__pe39__lane28_strm1_data_valid  ;

  output                                          pe39__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane29_strm0_data_mask   ;
  input                                           std__pe39__lane29_strm0_data_valid  ;

  output                                          pe39__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane29_strm1_data_mask   ;
  input                                           std__pe39__lane29_strm1_data_valid  ;

  output                                          pe39__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane30_strm0_data_mask   ;
  input                                           std__pe39__lane30_strm0_data_valid  ;

  output                                          pe39__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane30_strm1_data_mask   ;
  input                                           std__pe39__lane30_strm1_data_valid  ;

  output                                          pe39__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane31_strm0_data_mask   ;
  input                                           std__pe39__lane31_strm0_data_valid  ;

  output                                          pe39__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe39__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe39__lane31_strm1_data_mask   ;
  input                                           std__pe39__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe40__peId                ;
  input                                         sys__pe40__allSynchronized     ;
  output                                        pe40__sys__thisSynchronized    ;
  output                                        pe40__sys__ready               ;
  output                                        pe40__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe40__oob_cntl            ;
  input                                         std__pe40__oob_valid           ;
  output                                        pe40__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe40__oob_type            ;
  output                                          pe40__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane0_strm0_data_mask   ;
  input                                           std__pe40__lane0_strm0_data_valid  ;

  output                                          pe40__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane0_strm1_data_mask   ;
  input                                           std__pe40__lane0_strm1_data_valid  ;

  output                                          pe40__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane1_strm0_data_mask   ;
  input                                           std__pe40__lane1_strm0_data_valid  ;

  output                                          pe40__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane1_strm1_data_mask   ;
  input                                           std__pe40__lane1_strm1_data_valid  ;

  output                                          pe40__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane2_strm0_data_mask   ;
  input                                           std__pe40__lane2_strm0_data_valid  ;

  output                                          pe40__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane2_strm1_data_mask   ;
  input                                           std__pe40__lane2_strm1_data_valid  ;

  output                                          pe40__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane3_strm0_data_mask   ;
  input                                           std__pe40__lane3_strm0_data_valid  ;

  output                                          pe40__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane3_strm1_data_mask   ;
  input                                           std__pe40__lane3_strm1_data_valid  ;

  output                                          pe40__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane4_strm0_data_mask   ;
  input                                           std__pe40__lane4_strm0_data_valid  ;

  output                                          pe40__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane4_strm1_data_mask   ;
  input                                           std__pe40__lane4_strm1_data_valid  ;

  output                                          pe40__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane5_strm0_data_mask   ;
  input                                           std__pe40__lane5_strm0_data_valid  ;

  output                                          pe40__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane5_strm1_data_mask   ;
  input                                           std__pe40__lane5_strm1_data_valid  ;

  output                                          pe40__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane6_strm0_data_mask   ;
  input                                           std__pe40__lane6_strm0_data_valid  ;

  output                                          pe40__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane6_strm1_data_mask   ;
  input                                           std__pe40__lane6_strm1_data_valid  ;

  output                                          pe40__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane7_strm0_data_mask   ;
  input                                           std__pe40__lane7_strm0_data_valid  ;

  output                                          pe40__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane7_strm1_data_mask   ;
  input                                           std__pe40__lane7_strm1_data_valid  ;

  output                                          pe40__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane8_strm0_data_mask   ;
  input                                           std__pe40__lane8_strm0_data_valid  ;

  output                                          pe40__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane8_strm1_data_mask   ;
  input                                           std__pe40__lane8_strm1_data_valid  ;

  output                                          pe40__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane9_strm0_data_mask   ;
  input                                           std__pe40__lane9_strm0_data_valid  ;

  output                                          pe40__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane9_strm1_data_mask   ;
  input                                           std__pe40__lane9_strm1_data_valid  ;

  output                                          pe40__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane10_strm0_data_mask   ;
  input                                           std__pe40__lane10_strm0_data_valid  ;

  output                                          pe40__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane10_strm1_data_mask   ;
  input                                           std__pe40__lane10_strm1_data_valid  ;

  output                                          pe40__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane11_strm0_data_mask   ;
  input                                           std__pe40__lane11_strm0_data_valid  ;

  output                                          pe40__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane11_strm1_data_mask   ;
  input                                           std__pe40__lane11_strm1_data_valid  ;

  output                                          pe40__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane12_strm0_data_mask   ;
  input                                           std__pe40__lane12_strm0_data_valid  ;

  output                                          pe40__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane12_strm1_data_mask   ;
  input                                           std__pe40__lane12_strm1_data_valid  ;

  output                                          pe40__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane13_strm0_data_mask   ;
  input                                           std__pe40__lane13_strm0_data_valid  ;

  output                                          pe40__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane13_strm1_data_mask   ;
  input                                           std__pe40__lane13_strm1_data_valid  ;

  output                                          pe40__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane14_strm0_data_mask   ;
  input                                           std__pe40__lane14_strm0_data_valid  ;

  output                                          pe40__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane14_strm1_data_mask   ;
  input                                           std__pe40__lane14_strm1_data_valid  ;

  output                                          pe40__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane15_strm0_data_mask   ;
  input                                           std__pe40__lane15_strm0_data_valid  ;

  output                                          pe40__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane15_strm1_data_mask   ;
  input                                           std__pe40__lane15_strm1_data_valid  ;

  output                                          pe40__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane16_strm0_data_mask   ;
  input                                           std__pe40__lane16_strm0_data_valid  ;

  output                                          pe40__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane16_strm1_data_mask   ;
  input                                           std__pe40__lane16_strm1_data_valid  ;

  output                                          pe40__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane17_strm0_data_mask   ;
  input                                           std__pe40__lane17_strm0_data_valid  ;

  output                                          pe40__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane17_strm1_data_mask   ;
  input                                           std__pe40__lane17_strm1_data_valid  ;

  output                                          pe40__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane18_strm0_data_mask   ;
  input                                           std__pe40__lane18_strm0_data_valid  ;

  output                                          pe40__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane18_strm1_data_mask   ;
  input                                           std__pe40__lane18_strm1_data_valid  ;

  output                                          pe40__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane19_strm0_data_mask   ;
  input                                           std__pe40__lane19_strm0_data_valid  ;

  output                                          pe40__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane19_strm1_data_mask   ;
  input                                           std__pe40__lane19_strm1_data_valid  ;

  output                                          pe40__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane20_strm0_data_mask   ;
  input                                           std__pe40__lane20_strm0_data_valid  ;

  output                                          pe40__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane20_strm1_data_mask   ;
  input                                           std__pe40__lane20_strm1_data_valid  ;

  output                                          pe40__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane21_strm0_data_mask   ;
  input                                           std__pe40__lane21_strm0_data_valid  ;

  output                                          pe40__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane21_strm1_data_mask   ;
  input                                           std__pe40__lane21_strm1_data_valid  ;

  output                                          pe40__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane22_strm0_data_mask   ;
  input                                           std__pe40__lane22_strm0_data_valid  ;

  output                                          pe40__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane22_strm1_data_mask   ;
  input                                           std__pe40__lane22_strm1_data_valid  ;

  output                                          pe40__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane23_strm0_data_mask   ;
  input                                           std__pe40__lane23_strm0_data_valid  ;

  output                                          pe40__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane23_strm1_data_mask   ;
  input                                           std__pe40__lane23_strm1_data_valid  ;

  output                                          pe40__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane24_strm0_data_mask   ;
  input                                           std__pe40__lane24_strm0_data_valid  ;

  output                                          pe40__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane24_strm1_data_mask   ;
  input                                           std__pe40__lane24_strm1_data_valid  ;

  output                                          pe40__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane25_strm0_data_mask   ;
  input                                           std__pe40__lane25_strm0_data_valid  ;

  output                                          pe40__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane25_strm1_data_mask   ;
  input                                           std__pe40__lane25_strm1_data_valid  ;

  output                                          pe40__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane26_strm0_data_mask   ;
  input                                           std__pe40__lane26_strm0_data_valid  ;

  output                                          pe40__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane26_strm1_data_mask   ;
  input                                           std__pe40__lane26_strm1_data_valid  ;

  output                                          pe40__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane27_strm0_data_mask   ;
  input                                           std__pe40__lane27_strm0_data_valid  ;

  output                                          pe40__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane27_strm1_data_mask   ;
  input                                           std__pe40__lane27_strm1_data_valid  ;

  output                                          pe40__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane28_strm0_data_mask   ;
  input                                           std__pe40__lane28_strm0_data_valid  ;

  output                                          pe40__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane28_strm1_data_mask   ;
  input                                           std__pe40__lane28_strm1_data_valid  ;

  output                                          pe40__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane29_strm0_data_mask   ;
  input                                           std__pe40__lane29_strm0_data_valid  ;

  output                                          pe40__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane29_strm1_data_mask   ;
  input                                           std__pe40__lane29_strm1_data_valid  ;

  output                                          pe40__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane30_strm0_data_mask   ;
  input                                           std__pe40__lane30_strm0_data_valid  ;

  output                                          pe40__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane30_strm1_data_mask   ;
  input                                           std__pe40__lane30_strm1_data_valid  ;

  output                                          pe40__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane31_strm0_data_mask   ;
  input                                           std__pe40__lane31_strm0_data_valid  ;

  output                                          pe40__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe40__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe40__lane31_strm1_data_mask   ;
  input                                           std__pe40__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe41__peId                ;
  input                                         sys__pe41__allSynchronized     ;
  output                                        pe41__sys__thisSynchronized    ;
  output                                        pe41__sys__ready               ;
  output                                        pe41__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe41__oob_cntl            ;
  input                                         std__pe41__oob_valid           ;
  output                                        pe41__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe41__oob_type            ;
  output                                          pe41__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane0_strm0_data_mask   ;
  input                                           std__pe41__lane0_strm0_data_valid  ;

  output                                          pe41__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane0_strm1_data_mask   ;
  input                                           std__pe41__lane0_strm1_data_valid  ;

  output                                          pe41__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane1_strm0_data_mask   ;
  input                                           std__pe41__lane1_strm0_data_valid  ;

  output                                          pe41__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane1_strm1_data_mask   ;
  input                                           std__pe41__lane1_strm1_data_valid  ;

  output                                          pe41__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane2_strm0_data_mask   ;
  input                                           std__pe41__lane2_strm0_data_valid  ;

  output                                          pe41__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane2_strm1_data_mask   ;
  input                                           std__pe41__lane2_strm1_data_valid  ;

  output                                          pe41__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane3_strm0_data_mask   ;
  input                                           std__pe41__lane3_strm0_data_valid  ;

  output                                          pe41__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane3_strm1_data_mask   ;
  input                                           std__pe41__lane3_strm1_data_valid  ;

  output                                          pe41__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane4_strm0_data_mask   ;
  input                                           std__pe41__lane4_strm0_data_valid  ;

  output                                          pe41__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane4_strm1_data_mask   ;
  input                                           std__pe41__lane4_strm1_data_valid  ;

  output                                          pe41__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane5_strm0_data_mask   ;
  input                                           std__pe41__lane5_strm0_data_valid  ;

  output                                          pe41__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane5_strm1_data_mask   ;
  input                                           std__pe41__lane5_strm1_data_valid  ;

  output                                          pe41__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane6_strm0_data_mask   ;
  input                                           std__pe41__lane6_strm0_data_valid  ;

  output                                          pe41__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane6_strm1_data_mask   ;
  input                                           std__pe41__lane6_strm1_data_valid  ;

  output                                          pe41__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane7_strm0_data_mask   ;
  input                                           std__pe41__lane7_strm0_data_valid  ;

  output                                          pe41__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane7_strm1_data_mask   ;
  input                                           std__pe41__lane7_strm1_data_valid  ;

  output                                          pe41__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane8_strm0_data_mask   ;
  input                                           std__pe41__lane8_strm0_data_valid  ;

  output                                          pe41__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane8_strm1_data_mask   ;
  input                                           std__pe41__lane8_strm1_data_valid  ;

  output                                          pe41__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane9_strm0_data_mask   ;
  input                                           std__pe41__lane9_strm0_data_valid  ;

  output                                          pe41__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane9_strm1_data_mask   ;
  input                                           std__pe41__lane9_strm1_data_valid  ;

  output                                          pe41__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane10_strm0_data_mask   ;
  input                                           std__pe41__lane10_strm0_data_valid  ;

  output                                          pe41__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane10_strm1_data_mask   ;
  input                                           std__pe41__lane10_strm1_data_valid  ;

  output                                          pe41__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane11_strm0_data_mask   ;
  input                                           std__pe41__lane11_strm0_data_valid  ;

  output                                          pe41__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane11_strm1_data_mask   ;
  input                                           std__pe41__lane11_strm1_data_valid  ;

  output                                          pe41__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane12_strm0_data_mask   ;
  input                                           std__pe41__lane12_strm0_data_valid  ;

  output                                          pe41__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane12_strm1_data_mask   ;
  input                                           std__pe41__lane12_strm1_data_valid  ;

  output                                          pe41__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane13_strm0_data_mask   ;
  input                                           std__pe41__lane13_strm0_data_valid  ;

  output                                          pe41__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane13_strm1_data_mask   ;
  input                                           std__pe41__lane13_strm1_data_valid  ;

  output                                          pe41__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane14_strm0_data_mask   ;
  input                                           std__pe41__lane14_strm0_data_valid  ;

  output                                          pe41__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane14_strm1_data_mask   ;
  input                                           std__pe41__lane14_strm1_data_valid  ;

  output                                          pe41__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane15_strm0_data_mask   ;
  input                                           std__pe41__lane15_strm0_data_valid  ;

  output                                          pe41__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane15_strm1_data_mask   ;
  input                                           std__pe41__lane15_strm1_data_valid  ;

  output                                          pe41__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane16_strm0_data_mask   ;
  input                                           std__pe41__lane16_strm0_data_valid  ;

  output                                          pe41__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane16_strm1_data_mask   ;
  input                                           std__pe41__lane16_strm1_data_valid  ;

  output                                          pe41__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane17_strm0_data_mask   ;
  input                                           std__pe41__lane17_strm0_data_valid  ;

  output                                          pe41__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane17_strm1_data_mask   ;
  input                                           std__pe41__lane17_strm1_data_valid  ;

  output                                          pe41__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane18_strm0_data_mask   ;
  input                                           std__pe41__lane18_strm0_data_valid  ;

  output                                          pe41__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane18_strm1_data_mask   ;
  input                                           std__pe41__lane18_strm1_data_valid  ;

  output                                          pe41__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane19_strm0_data_mask   ;
  input                                           std__pe41__lane19_strm0_data_valid  ;

  output                                          pe41__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane19_strm1_data_mask   ;
  input                                           std__pe41__lane19_strm1_data_valid  ;

  output                                          pe41__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane20_strm0_data_mask   ;
  input                                           std__pe41__lane20_strm0_data_valid  ;

  output                                          pe41__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane20_strm1_data_mask   ;
  input                                           std__pe41__lane20_strm1_data_valid  ;

  output                                          pe41__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane21_strm0_data_mask   ;
  input                                           std__pe41__lane21_strm0_data_valid  ;

  output                                          pe41__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane21_strm1_data_mask   ;
  input                                           std__pe41__lane21_strm1_data_valid  ;

  output                                          pe41__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane22_strm0_data_mask   ;
  input                                           std__pe41__lane22_strm0_data_valid  ;

  output                                          pe41__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane22_strm1_data_mask   ;
  input                                           std__pe41__lane22_strm1_data_valid  ;

  output                                          pe41__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane23_strm0_data_mask   ;
  input                                           std__pe41__lane23_strm0_data_valid  ;

  output                                          pe41__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane23_strm1_data_mask   ;
  input                                           std__pe41__lane23_strm1_data_valid  ;

  output                                          pe41__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane24_strm0_data_mask   ;
  input                                           std__pe41__lane24_strm0_data_valid  ;

  output                                          pe41__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane24_strm1_data_mask   ;
  input                                           std__pe41__lane24_strm1_data_valid  ;

  output                                          pe41__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane25_strm0_data_mask   ;
  input                                           std__pe41__lane25_strm0_data_valid  ;

  output                                          pe41__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane25_strm1_data_mask   ;
  input                                           std__pe41__lane25_strm1_data_valid  ;

  output                                          pe41__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane26_strm0_data_mask   ;
  input                                           std__pe41__lane26_strm0_data_valid  ;

  output                                          pe41__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane26_strm1_data_mask   ;
  input                                           std__pe41__lane26_strm1_data_valid  ;

  output                                          pe41__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane27_strm0_data_mask   ;
  input                                           std__pe41__lane27_strm0_data_valid  ;

  output                                          pe41__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane27_strm1_data_mask   ;
  input                                           std__pe41__lane27_strm1_data_valid  ;

  output                                          pe41__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane28_strm0_data_mask   ;
  input                                           std__pe41__lane28_strm0_data_valid  ;

  output                                          pe41__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane28_strm1_data_mask   ;
  input                                           std__pe41__lane28_strm1_data_valid  ;

  output                                          pe41__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane29_strm0_data_mask   ;
  input                                           std__pe41__lane29_strm0_data_valid  ;

  output                                          pe41__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane29_strm1_data_mask   ;
  input                                           std__pe41__lane29_strm1_data_valid  ;

  output                                          pe41__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane30_strm0_data_mask   ;
  input                                           std__pe41__lane30_strm0_data_valid  ;

  output                                          pe41__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane30_strm1_data_mask   ;
  input                                           std__pe41__lane30_strm1_data_valid  ;

  output                                          pe41__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane31_strm0_data_mask   ;
  input                                           std__pe41__lane31_strm0_data_valid  ;

  output                                          pe41__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe41__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe41__lane31_strm1_data_mask   ;
  input                                           std__pe41__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe42__peId                ;
  input                                         sys__pe42__allSynchronized     ;
  output                                        pe42__sys__thisSynchronized    ;
  output                                        pe42__sys__ready               ;
  output                                        pe42__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe42__oob_cntl            ;
  input                                         std__pe42__oob_valid           ;
  output                                        pe42__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe42__oob_type            ;
  output                                          pe42__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane0_strm0_data_mask   ;
  input                                           std__pe42__lane0_strm0_data_valid  ;

  output                                          pe42__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane0_strm1_data_mask   ;
  input                                           std__pe42__lane0_strm1_data_valid  ;

  output                                          pe42__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane1_strm0_data_mask   ;
  input                                           std__pe42__lane1_strm0_data_valid  ;

  output                                          pe42__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane1_strm1_data_mask   ;
  input                                           std__pe42__lane1_strm1_data_valid  ;

  output                                          pe42__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane2_strm0_data_mask   ;
  input                                           std__pe42__lane2_strm0_data_valid  ;

  output                                          pe42__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane2_strm1_data_mask   ;
  input                                           std__pe42__lane2_strm1_data_valid  ;

  output                                          pe42__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane3_strm0_data_mask   ;
  input                                           std__pe42__lane3_strm0_data_valid  ;

  output                                          pe42__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane3_strm1_data_mask   ;
  input                                           std__pe42__lane3_strm1_data_valid  ;

  output                                          pe42__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane4_strm0_data_mask   ;
  input                                           std__pe42__lane4_strm0_data_valid  ;

  output                                          pe42__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane4_strm1_data_mask   ;
  input                                           std__pe42__lane4_strm1_data_valid  ;

  output                                          pe42__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane5_strm0_data_mask   ;
  input                                           std__pe42__lane5_strm0_data_valid  ;

  output                                          pe42__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane5_strm1_data_mask   ;
  input                                           std__pe42__lane5_strm1_data_valid  ;

  output                                          pe42__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane6_strm0_data_mask   ;
  input                                           std__pe42__lane6_strm0_data_valid  ;

  output                                          pe42__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane6_strm1_data_mask   ;
  input                                           std__pe42__lane6_strm1_data_valid  ;

  output                                          pe42__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane7_strm0_data_mask   ;
  input                                           std__pe42__lane7_strm0_data_valid  ;

  output                                          pe42__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane7_strm1_data_mask   ;
  input                                           std__pe42__lane7_strm1_data_valid  ;

  output                                          pe42__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane8_strm0_data_mask   ;
  input                                           std__pe42__lane8_strm0_data_valid  ;

  output                                          pe42__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane8_strm1_data_mask   ;
  input                                           std__pe42__lane8_strm1_data_valid  ;

  output                                          pe42__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane9_strm0_data_mask   ;
  input                                           std__pe42__lane9_strm0_data_valid  ;

  output                                          pe42__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane9_strm1_data_mask   ;
  input                                           std__pe42__lane9_strm1_data_valid  ;

  output                                          pe42__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane10_strm0_data_mask   ;
  input                                           std__pe42__lane10_strm0_data_valid  ;

  output                                          pe42__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane10_strm1_data_mask   ;
  input                                           std__pe42__lane10_strm1_data_valid  ;

  output                                          pe42__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane11_strm0_data_mask   ;
  input                                           std__pe42__lane11_strm0_data_valid  ;

  output                                          pe42__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane11_strm1_data_mask   ;
  input                                           std__pe42__lane11_strm1_data_valid  ;

  output                                          pe42__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane12_strm0_data_mask   ;
  input                                           std__pe42__lane12_strm0_data_valid  ;

  output                                          pe42__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane12_strm1_data_mask   ;
  input                                           std__pe42__lane12_strm1_data_valid  ;

  output                                          pe42__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane13_strm0_data_mask   ;
  input                                           std__pe42__lane13_strm0_data_valid  ;

  output                                          pe42__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane13_strm1_data_mask   ;
  input                                           std__pe42__lane13_strm1_data_valid  ;

  output                                          pe42__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane14_strm0_data_mask   ;
  input                                           std__pe42__lane14_strm0_data_valid  ;

  output                                          pe42__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane14_strm1_data_mask   ;
  input                                           std__pe42__lane14_strm1_data_valid  ;

  output                                          pe42__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane15_strm0_data_mask   ;
  input                                           std__pe42__lane15_strm0_data_valid  ;

  output                                          pe42__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane15_strm1_data_mask   ;
  input                                           std__pe42__lane15_strm1_data_valid  ;

  output                                          pe42__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane16_strm0_data_mask   ;
  input                                           std__pe42__lane16_strm0_data_valid  ;

  output                                          pe42__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane16_strm1_data_mask   ;
  input                                           std__pe42__lane16_strm1_data_valid  ;

  output                                          pe42__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane17_strm0_data_mask   ;
  input                                           std__pe42__lane17_strm0_data_valid  ;

  output                                          pe42__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane17_strm1_data_mask   ;
  input                                           std__pe42__lane17_strm1_data_valid  ;

  output                                          pe42__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane18_strm0_data_mask   ;
  input                                           std__pe42__lane18_strm0_data_valid  ;

  output                                          pe42__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane18_strm1_data_mask   ;
  input                                           std__pe42__lane18_strm1_data_valid  ;

  output                                          pe42__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane19_strm0_data_mask   ;
  input                                           std__pe42__lane19_strm0_data_valid  ;

  output                                          pe42__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane19_strm1_data_mask   ;
  input                                           std__pe42__lane19_strm1_data_valid  ;

  output                                          pe42__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane20_strm0_data_mask   ;
  input                                           std__pe42__lane20_strm0_data_valid  ;

  output                                          pe42__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane20_strm1_data_mask   ;
  input                                           std__pe42__lane20_strm1_data_valid  ;

  output                                          pe42__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane21_strm0_data_mask   ;
  input                                           std__pe42__lane21_strm0_data_valid  ;

  output                                          pe42__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane21_strm1_data_mask   ;
  input                                           std__pe42__lane21_strm1_data_valid  ;

  output                                          pe42__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane22_strm0_data_mask   ;
  input                                           std__pe42__lane22_strm0_data_valid  ;

  output                                          pe42__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane22_strm1_data_mask   ;
  input                                           std__pe42__lane22_strm1_data_valid  ;

  output                                          pe42__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane23_strm0_data_mask   ;
  input                                           std__pe42__lane23_strm0_data_valid  ;

  output                                          pe42__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane23_strm1_data_mask   ;
  input                                           std__pe42__lane23_strm1_data_valid  ;

  output                                          pe42__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane24_strm0_data_mask   ;
  input                                           std__pe42__lane24_strm0_data_valid  ;

  output                                          pe42__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane24_strm1_data_mask   ;
  input                                           std__pe42__lane24_strm1_data_valid  ;

  output                                          pe42__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane25_strm0_data_mask   ;
  input                                           std__pe42__lane25_strm0_data_valid  ;

  output                                          pe42__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane25_strm1_data_mask   ;
  input                                           std__pe42__lane25_strm1_data_valid  ;

  output                                          pe42__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane26_strm0_data_mask   ;
  input                                           std__pe42__lane26_strm0_data_valid  ;

  output                                          pe42__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane26_strm1_data_mask   ;
  input                                           std__pe42__lane26_strm1_data_valid  ;

  output                                          pe42__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane27_strm0_data_mask   ;
  input                                           std__pe42__lane27_strm0_data_valid  ;

  output                                          pe42__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane27_strm1_data_mask   ;
  input                                           std__pe42__lane27_strm1_data_valid  ;

  output                                          pe42__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane28_strm0_data_mask   ;
  input                                           std__pe42__lane28_strm0_data_valid  ;

  output                                          pe42__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane28_strm1_data_mask   ;
  input                                           std__pe42__lane28_strm1_data_valid  ;

  output                                          pe42__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane29_strm0_data_mask   ;
  input                                           std__pe42__lane29_strm0_data_valid  ;

  output                                          pe42__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane29_strm1_data_mask   ;
  input                                           std__pe42__lane29_strm1_data_valid  ;

  output                                          pe42__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane30_strm0_data_mask   ;
  input                                           std__pe42__lane30_strm0_data_valid  ;

  output                                          pe42__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane30_strm1_data_mask   ;
  input                                           std__pe42__lane30_strm1_data_valid  ;

  output                                          pe42__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane31_strm0_data_mask   ;
  input                                           std__pe42__lane31_strm0_data_valid  ;

  output                                          pe42__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe42__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe42__lane31_strm1_data_mask   ;
  input                                           std__pe42__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe43__peId                ;
  input                                         sys__pe43__allSynchronized     ;
  output                                        pe43__sys__thisSynchronized    ;
  output                                        pe43__sys__ready               ;
  output                                        pe43__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe43__oob_cntl            ;
  input                                         std__pe43__oob_valid           ;
  output                                        pe43__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe43__oob_type            ;
  output                                          pe43__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane0_strm0_data_mask   ;
  input                                           std__pe43__lane0_strm0_data_valid  ;

  output                                          pe43__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane0_strm1_data_mask   ;
  input                                           std__pe43__lane0_strm1_data_valid  ;

  output                                          pe43__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane1_strm0_data_mask   ;
  input                                           std__pe43__lane1_strm0_data_valid  ;

  output                                          pe43__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane1_strm1_data_mask   ;
  input                                           std__pe43__lane1_strm1_data_valid  ;

  output                                          pe43__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane2_strm0_data_mask   ;
  input                                           std__pe43__lane2_strm0_data_valid  ;

  output                                          pe43__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane2_strm1_data_mask   ;
  input                                           std__pe43__lane2_strm1_data_valid  ;

  output                                          pe43__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane3_strm0_data_mask   ;
  input                                           std__pe43__lane3_strm0_data_valid  ;

  output                                          pe43__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane3_strm1_data_mask   ;
  input                                           std__pe43__lane3_strm1_data_valid  ;

  output                                          pe43__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane4_strm0_data_mask   ;
  input                                           std__pe43__lane4_strm0_data_valid  ;

  output                                          pe43__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane4_strm1_data_mask   ;
  input                                           std__pe43__lane4_strm1_data_valid  ;

  output                                          pe43__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane5_strm0_data_mask   ;
  input                                           std__pe43__lane5_strm0_data_valid  ;

  output                                          pe43__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane5_strm1_data_mask   ;
  input                                           std__pe43__lane5_strm1_data_valid  ;

  output                                          pe43__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane6_strm0_data_mask   ;
  input                                           std__pe43__lane6_strm0_data_valid  ;

  output                                          pe43__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane6_strm1_data_mask   ;
  input                                           std__pe43__lane6_strm1_data_valid  ;

  output                                          pe43__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane7_strm0_data_mask   ;
  input                                           std__pe43__lane7_strm0_data_valid  ;

  output                                          pe43__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane7_strm1_data_mask   ;
  input                                           std__pe43__lane7_strm1_data_valid  ;

  output                                          pe43__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane8_strm0_data_mask   ;
  input                                           std__pe43__lane8_strm0_data_valid  ;

  output                                          pe43__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane8_strm1_data_mask   ;
  input                                           std__pe43__lane8_strm1_data_valid  ;

  output                                          pe43__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane9_strm0_data_mask   ;
  input                                           std__pe43__lane9_strm0_data_valid  ;

  output                                          pe43__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane9_strm1_data_mask   ;
  input                                           std__pe43__lane9_strm1_data_valid  ;

  output                                          pe43__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane10_strm0_data_mask   ;
  input                                           std__pe43__lane10_strm0_data_valid  ;

  output                                          pe43__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane10_strm1_data_mask   ;
  input                                           std__pe43__lane10_strm1_data_valid  ;

  output                                          pe43__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane11_strm0_data_mask   ;
  input                                           std__pe43__lane11_strm0_data_valid  ;

  output                                          pe43__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane11_strm1_data_mask   ;
  input                                           std__pe43__lane11_strm1_data_valid  ;

  output                                          pe43__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane12_strm0_data_mask   ;
  input                                           std__pe43__lane12_strm0_data_valid  ;

  output                                          pe43__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane12_strm1_data_mask   ;
  input                                           std__pe43__lane12_strm1_data_valid  ;

  output                                          pe43__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane13_strm0_data_mask   ;
  input                                           std__pe43__lane13_strm0_data_valid  ;

  output                                          pe43__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane13_strm1_data_mask   ;
  input                                           std__pe43__lane13_strm1_data_valid  ;

  output                                          pe43__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane14_strm0_data_mask   ;
  input                                           std__pe43__lane14_strm0_data_valid  ;

  output                                          pe43__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane14_strm1_data_mask   ;
  input                                           std__pe43__lane14_strm1_data_valid  ;

  output                                          pe43__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane15_strm0_data_mask   ;
  input                                           std__pe43__lane15_strm0_data_valid  ;

  output                                          pe43__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane15_strm1_data_mask   ;
  input                                           std__pe43__lane15_strm1_data_valid  ;

  output                                          pe43__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane16_strm0_data_mask   ;
  input                                           std__pe43__lane16_strm0_data_valid  ;

  output                                          pe43__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane16_strm1_data_mask   ;
  input                                           std__pe43__lane16_strm1_data_valid  ;

  output                                          pe43__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane17_strm0_data_mask   ;
  input                                           std__pe43__lane17_strm0_data_valid  ;

  output                                          pe43__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane17_strm1_data_mask   ;
  input                                           std__pe43__lane17_strm1_data_valid  ;

  output                                          pe43__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane18_strm0_data_mask   ;
  input                                           std__pe43__lane18_strm0_data_valid  ;

  output                                          pe43__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane18_strm1_data_mask   ;
  input                                           std__pe43__lane18_strm1_data_valid  ;

  output                                          pe43__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane19_strm0_data_mask   ;
  input                                           std__pe43__lane19_strm0_data_valid  ;

  output                                          pe43__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane19_strm1_data_mask   ;
  input                                           std__pe43__lane19_strm1_data_valid  ;

  output                                          pe43__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane20_strm0_data_mask   ;
  input                                           std__pe43__lane20_strm0_data_valid  ;

  output                                          pe43__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane20_strm1_data_mask   ;
  input                                           std__pe43__lane20_strm1_data_valid  ;

  output                                          pe43__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane21_strm0_data_mask   ;
  input                                           std__pe43__lane21_strm0_data_valid  ;

  output                                          pe43__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane21_strm1_data_mask   ;
  input                                           std__pe43__lane21_strm1_data_valid  ;

  output                                          pe43__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane22_strm0_data_mask   ;
  input                                           std__pe43__lane22_strm0_data_valid  ;

  output                                          pe43__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane22_strm1_data_mask   ;
  input                                           std__pe43__lane22_strm1_data_valid  ;

  output                                          pe43__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane23_strm0_data_mask   ;
  input                                           std__pe43__lane23_strm0_data_valid  ;

  output                                          pe43__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane23_strm1_data_mask   ;
  input                                           std__pe43__lane23_strm1_data_valid  ;

  output                                          pe43__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane24_strm0_data_mask   ;
  input                                           std__pe43__lane24_strm0_data_valid  ;

  output                                          pe43__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane24_strm1_data_mask   ;
  input                                           std__pe43__lane24_strm1_data_valid  ;

  output                                          pe43__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane25_strm0_data_mask   ;
  input                                           std__pe43__lane25_strm0_data_valid  ;

  output                                          pe43__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane25_strm1_data_mask   ;
  input                                           std__pe43__lane25_strm1_data_valid  ;

  output                                          pe43__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane26_strm0_data_mask   ;
  input                                           std__pe43__lane26_strm0_data_valid  ;

  output                                          pe43__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane26_strm1_data_mask   ;
  input                                           std__pe43__lane26_strm1_data_valid  ;

  output                                          pe43__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane27_strm0_data_mask   ;
  input                                           std__pe43__lane27_strm0_data_valid  ;

  output                                          pe43__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane27_strm1_data_mask   ;
  input                                           std__pe43__lane27_strm1_data_valid  ;

  output                                          pe43__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane28_strm0_data_mask   ;
  input                                           std__pe43__lane28_strm0_data_valid  ;

  output                                          pe43__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane28_strm1_data_mask   ;
  input                                           std__pe43__lane28_strm1_data_valid  ;

  output                                          pe43__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane29_strm0_data_mask   ;
  input                                           std__pe43__lane29_strm0_data_valid  ;

  output                                          pe43__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane29_strm1_data_mask   ;
  input                                           std__pe43__lane29_strm1_data_valid  ;

  output                                          pe43__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane30_strm0_data_mask   ;
  input                                           std__pe43__lane30_strm0_data_valid  ;

  output                                          pe43__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane30_strm1_data_mask   ;
  input                                           std__pe43__lane30_strm1_data_valid  ;

  output                                          pe43__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane31_strm0_data_mask   ;
  input                                           std__pe43__lane31_strm0_data_valid  ;

  output                                          pe43__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe43__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe43__lane31_strm1_data_mask   ;
  input                                           std__pe43__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe44__peId                ;
  input                                         sys__pe44__allSynchronized     ;
  output                                        pe44__sys__thisSynchronized    ;
  output                                        pe44__sys__ready               ;
  output                                        pe44__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe44__oob_cntl            ;
  input                                         std__pe44__oob_valid           ;
  output                                        pe44__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe44__oob_type            ;
  output                                          pe44__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane0_strm0_data_mask   ;
  input                                           std__pe44__lane0_strm0_data_valid  ;

  output                                          pe44__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane0_strm1_data_mask   ;
  input                                           std__pe44__lane0_strm1_data_valid  ;

  output                                          pe44__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane1_strm0_data_mask   ;
  input                                           std__pe44__lane1_strm0_data_valid  ;

  output                                          pe44__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane1_strm1_data_mask   ;
  input                                           std__pe44__lane1_strm1_data_valid  ;

  output                                          pe44__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane2_strm0_data_mask   ;
  input                                           std__pe44__lane2_strm0_data_valid  ;

  output                                          pe44__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane2_strm1_data_mask   ;
  input                                           std__pe44__lane2_strm1_data_valid  ;

  output                                          pe44__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane3_strm0_data_mask   ;
  input                                           std__pe44__lane3_strm0_data_valid  ;

  output                                          pe44__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane3_strm1_data_mask   ;
  input                                           std__pe44__lane3_strm1_data_valid  ;

  output                                          pe44__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane4_strm0_data_mask   ;
  input                                           std__pe44__lane4_strm0_data_valid  ;

  output                                          pe44__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane4_strm1_data_mask   ;
  input                                           std__pe44__lane4_strm1_data_valid  ;

  output                                          pe44__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane5_strm0_data_mask   ;
  input                                           std__pe44__lane5_strm0_data_valid  ;

  output                                          pe44__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane5_strm1_data_mask   ;
  input                                           std__pe44__lane5_strm1_data_valid  ;

  output                                          pe44__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane6_strm0_data_mask   ;
  input                                           std__pe44__lane6_strm0_data_valid  ;

  output                                          pe44__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane6_strm1_data_mask   ;
  input                                           std__pe44__lane6_strm1_data_valid  ;

  output                                          pe44__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane7_strm0_data_mask   ;
  input                                           std__pe44__lane7_strm0_data_valid  ;

  output                                          pe44__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane7_strm1_data_mask   ;
  input                                           std__pe44__lane7_strm1_data_valid  ;

  output                                          pe44__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane8_strm0_data_mask   ;
  input                                           std__pe44__lane8_strm0_data_valid  ;

  output                                          pe44__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane8_strm1_data_mask   ;
  input                                           std__pe44__lane8_strm1_data_valid  ;

  output                                          pe44__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane9_strm0_data_mask   ;
  input                                           std__pe44__lane9_strm0_data_valid  ;

  output                                          pe44__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane9_strm1_data_mask   ;
  input                                           std__pe44__lane9_strm1_data_valid  ;

  output                                          pe44__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane10_strm0_data_mask   ;
  input                                           std__pe44__lane10_strm0_data_valid  ;

  output                                          pe44__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane10_strm1_data_mask   ;
  input                                           std__pe44__lane10_strm1_data_valid  ;

  output                                          pe44__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane11_strm0_data_mask   ;
  input                                           std__pe44__lane11_strm0_data_valid  ;

  output                                          pe44__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane11_strm1_data_mask   ;
  input                                           std__pe44__lane11_strm1_data_valid  ;

  output                                          pe44__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane12_strm0_data_mask   ;
  input                                           std__pe44__lane12_strm0_data_valid  ;

  output                                          pe44__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane12_strm1_data_mask   ;
  input                                           std__pe44__lane12_strm1_data_valid  ;

  output                                          pe44__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane13_strm0_data_mask   ;
  input                                           std__pe44__lane13_strm0_data_valid  ;

  output                                          pe44__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane13_strm1_data_mask   ;
  input                                           std__pe44__lane13_strm1_data_valid  ;

  output                                          pe44__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane14_strm0_data_mask   ;
  input                                           std__pe44__lane14_strm0_data_valid  ;

  output                                          pe44__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane14_strm1_data_mask   ;
  input                                           std__pe44__lane14_strm1_data_valid  ;

  output                                          pe44__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane15_strm0_data_mask   ;
  input                                           std__pe44__lane15_strm0_data_valid  ;

  output                                          pe44__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane15_strm1_data_mask   ;
  input                                           std__pe44__lane15_strm1_data_valid  ;

  output                                          pe44__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane16_strm0_data_mask   ;
  input                                           std__pe44__lane16_strm0_data_valid  ;

  output                                          pe44__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane16_strm1_data_mask   ;
  input                                           std__pe44__lane16_strm1_data_valid  ;

  output                                          pe44__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane17_strm0_data_mask   ;
  input                                           std__pe44__lane17_strm0_data_valid  ;

  output                                          pe44__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane17_strm1_data_mask   ;
  input                                           std__pe44__lane17_strm1_data_valid  ;

  output                                          pe44__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane18_strm0_data_mask   ;
  input                                           std__pe44__lane18_strm0_data_valid  ;

  output                                          pe44__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane18_strm1_data_mask   ;
  input                                           std__pe44__lane18_strm1_data_valid  ;

  output                                          pe44__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane19_strm0_data_mask   ;
  input                                           std__pe44__lane19_strm0_data_valid  ;

  output                                          pe44__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane19_strm1_data_mask   ;
  input                                           std__pe44__lane19_strm1_data_valid  ;

  output                                          pe44__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane20_strm0_data_mask   ;
  input                                           std__pe44__lane20_strm0_data_valid  ;

  output                                          pe44__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane20_strm1_data_mask   ;
  input                                           std__pe44__lane20_strm1_data_valid  ;

  output                                          pe44__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane21_strm0_data_mask   ;
  input                                           std__pe44__lane21_strm0_data_valid  ;

  output                                          pe44__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane21_strm1_data_mask   ;
  input                                           std__pe44__lane21_strm1_data_valid  ;

  output                                          pe44__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane22_strm0_data_mask   ;
  input                                           std__pe44__lane22_strm0_data_valid  ;

  output                                          pe44__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane22_strm1_data_mask   ;
  input                                           std__pe44__lane22_strm1_data_valid  ;

  output                                          pe44__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane23_strm0_data_mask   ;
  input                                           std__pe44__lane23_strm0_data_valid  ;

  output                                          pe44__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane23_strm1_data_mask   ;
  input                                           std__pe44__lane23_strm1_data_valid  ;

  output                                          pe44__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane24_strm0_data_mask   ;
  input                                           std__pe44__lane24_strm0_data_valid  ;

  output                                          pe44__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane24_strm1_data_mask   ;
  input                                           std__pe44__lane24_strm1_data_valid  ;

  output                                          pe44__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane25_strm0_data_mask   ;
  input                                           std__pe44__lane25_strm0_data_valid  ;

  output                                          pe44__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane25_strm1_data_mask   ;
  input                                           std__pe44__lane25_strm1_data_valid  ;

  output                                          pe44__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane26_strm0_data_mask   ;
  input                                           std__pe44__lane26_strm0_data_valid  ;

  output                                          pe44__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane26_strm1_data_mask   ;
  input                                           std__pe44__lane26_strm1_data_valid  ;

  output                                          pe44__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane27_strm0_data_mask   ;
  input                                           std__pe44__lane27_strm0_data_valid  ;

  output                                          pe44__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane27_strm1_data_mask   ;
  input                                           std__pe44__lane27_strm1_data_valid  ;

  output                                          pe44__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane28_strm0_data_mask   ;
  input                                           std__pe44__lane28_strm0_data_valid  ;

  output                                          pe44__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane28_strm1_data_mask   ;
  input                                           std__pe44__lane28_strm1_data_valid  ;

  output                                          pe44__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane29_strm0_data_mask   ;
  input                                           std__pe44__lane29_strm0_data_valid  ;

  output                                          pe44__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane29_strm1_data_mask   ;
  input                                           std__pe44__lane29_strm1_data_valid  ;

  output                                          pe44__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane30_strm0_data_mask   ;
  input                                           std__pe44__lane30_strm0_data_valid  ;

  output                                          pe44__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane30_strm1_data_mask   ;
  input                                           std__pe44__lane30_strm1_data_valid  ;

  output                                          pe44__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane31_strm0_data_mask   ;
  input                                           std__pe44__lane31_strm0_data_valid  ;

  output                                          pe44__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe44__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe44__lane31_strm1_data_mask   ;
  input                                           std__pe44__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe45__peId                ;
  input                                         sys__pe45__allSynchronized     ;
  output                                        pe45__sys__thisSynchronized    ;
  output                                        pe45__sys__ready               ;
  output                                        pe45__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe45__oob_cntl            ;
  input                                         std__pe45__oob_valid           ;
  output                                        pe45__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe45__oob_type            ;
  output                                          pe45__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane0_strm0_data_mask   ;
  input                                           std__pe45__lane0_strm0_data_valid  ;

  output                                          pe45__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane0_strm1_data_mask   ;
  input                                           std__pe45__lane0_strm1_data_valid  ;

  output                                          pe45__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane1_strm0_data_mask   ;
  input                                           std__pe45__lane1_strm0_data_valid  ;

  output                                          pe45__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane1_strm1_data_mask   ;
  input                                           std__pe45__lane1_strm1_data_valid  ;

  output                                          pe45__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane2_strm0_data_mask   ;
  input                                           std__pe45__lane2_strm0_data_valid  ;

  output                                          pe45__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane2_strm1_data_mask   ;
  input                                           std__pe45__lane2_strm1_data_valid  ;

  output                                          pe45__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane3_strm0_data_mask   ;
  input                                           std__pe45__lane3_strm0_data_valid  ;

  output                                          pe45__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane3_strm1_data_mask   ;
  input                                           std__pe45__lane3_strm1_data_valid  ;

  output                                          pe45__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane4_strm0_data_mask   ;
  input                                           std__pe45__lane4_strm0_data_valid  ;

  output                                          pe45__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane4_strm1_data_mask   ;
  input                                           std__pe45__lane4_strm1_data_valid  ;

  output                                          pe45__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane5_strm0_data_mask   ;
  input                                           std__pe45__lane5_strm0_data_valid  ;

  output                                          pe45__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane5_strm1_data_mask   ;
  input                                           std__pe45__lane5_strm1_data_valid  ;

  output                                          pe45__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane6_strm0_data_mask   ;
  input                                           std__pe45__lane6_strm0_data_valid  ;

  output                                          pe45__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane6_strm1_data_mask   ;
  input                                           std__pe45__lane6_strm1_data_valid  ;

  output                                          pe45__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane7_strm0_data_mask   ;
  input                                           std__pe45__lane7_strm0_data_valid  ;

  output                                          pe45__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane7_strm1_data_mask   ;
  input                                           std__pe45__lane7_strm1_data_valid  ;

  output                                          pe45__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane8_strm0_data_mask   ;
  input                                           std__pe45__lane8_strm0_data_valid  ;

  output                                          pe45__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane8_strm1_data_mask   ;
  input                                           std__pe45__lane8_strm1_data_valid  ;

  output                                          pe45__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane9_strm0_data_mask   ;
  input                                           std__pe45__lane9_strm0_data_valid  ;

  output                                          pe45__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane9_strm1_data_mask   ;
  input                                           std__pe45__lane9_strm1_data_valid  ;

  output                                          pe45__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane10_strm0_data_mask   ;
  input                                           std__pe45__lane10_strm0_data_valid  ;

  output                                          pe45__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane10_strm1_data_mask   ;
  input                                           std__pe45__lane10_strm1_data_valid  ;

  output                                          pe45__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane11_strm0_data_mask   ;
  input                                           std__pe45__lane11_strm0_data_valid  ;

  output                                          pe45__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane11_strm1_data_mask   ;
  input                                           std__pe45__lane11_strm1_data_valid  ;

  output                                          pe45__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane12_strm0_data_mask   ;
  input                                           std__pe45__lane12_strm0_data_valid  ;

  output                                          pe45__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane12_strm1_data_mask   ;
  input                                           std__pe45__lane12_strm1_data_valid  ;

  output                                          pe45__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane13_strm0_data_mask   ;
  input                                           std__pe45__lane13_strm0_data_valid  ;

  output                                          pe45__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane13_strm1_data_mask   ;
  input                                           std__pe45__lane13_strm1_data_valid  ;

  output                                          pe45__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane14_strm0_data_mask   ;
  input                                           std__pe45__lane14_strm0_data_valid  ;

  output                                          pe45__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane14_strm1_data_mask   ;
  input                                           std__pe45__lane14_strm1_data_valid  ;

  output                                          pe45__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane15_strm0_data_mask   ;
  input                                           std__pe45__lane15_strm0_data_valid  ;

  output                                          pe45__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane15_strm1_data_mask   ;
  input                                           std__pe45__lane15_strm1_data_valid  ;

  output                                          pe45__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane16_strm0_data_mask   ;
  input                                           std__pe45__lane16_strm0_data_valid  ;

  output                                          pe45__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane16_strm1_data_mask   ;
  input                                           std__pe45__lane16_strm1_data_valid  ;

  output                                          pe45__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane17_strm0_data_mask   ;
  input                                           std__pe45__lane17_strm0_data_valid  ;

  output                                          pe45__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane17_strm1_data_mask   ;
  input                                           std__pe45__lane17_strm1_data_valid  ;

  output                                          pe45__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane18_strm0_data_mask   ;
  input                                           std__pe45__lane18_strm0_data_valid  ;

  output                                          pe45__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane18_strm1_data_mask   ;
  input                                           std__pe45__lane18_strm1_data_valid  ;

  output                                          pe45__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane19_strm0_data_mask   ;
  input                                           std__pe45__lane19_strm0_data_valid  ;

  output                                          pe45__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane19_strm1_data_mask   ;
  input                                           std__pe45__lane19_strm1_data_valid  ;

  output                                          pe45__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane20_strm0_data_mask   ;
  input                                           std__pe45__lane20_strm0_data_valid  ;

  output                                          pe45__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane20_strm1_data_mask   ;
  input                                           std__pe45__lane20_strm1_data_valid  ;

  output                                          pe45__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane21_strm0_data_mask   ;
  input                                           std__pe45__lane21_strm0_data_valid  ;

  output                                          pe45__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane21_strm1_data_mask   ;
  input                                           std__pe45__lane21_strm1_data_valid  ;

  output                                          pe45__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane22_strm0_data_mask   ;
  input                                           std__pe45__lane22_strm0_data_valid  ;

  output                                          pe45__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane22_strm1_data_mask   ;
  input                                           std__pe45__lane22_strm1_data_valid  ;

  output                                          pe45__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane23_strm0_data_mask   ;
  input                                           std__pe45__lane23_strm0_data_valid  ;

  output                                          pe45__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane23_strm1_data_mask   ;
  input                                           std__pe45__lane23_strm1_data_valid  ;

  output                                          pe45__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane24_strm0_data_mask   ;
  input                                           std__pe45__lane24_strm0_data_valid  ;

  output                                          pe45__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane24_strm1_data_mask   ;
  input                                           std__pe45__lane24_strm1_data_valid  ;

  output                                          pe45__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane25_strm0_data_mask   ;
  input                                           std__pe45__lane25_strm0_data_valid  ;

  output                                          pe45__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane25_strm1_data_mask   ;
  input                                           std__pe45__lane25_strm1_data_valid  ;

  output                                          pe45__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane26_strm0_data_mask   ;
  input                                           std__pe45__lane26_strm0_data_valid  ;

  output                                          pe45__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane26_strm1_data_mask   ;
  input                                           std__pe45__lane26_strm1_data_valid  ;

  output                                          pe45__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane27_strm0_data_mask   ;
  input                                           std__pe45__lane27_strm0_data_valid  ;

  output                                          pe45__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane27_strm1_data_mask   ;
  input                                           std__pe45__lane27_strm1_data_valid  ;

  output                                          pe45__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane28_strm0_data_mask   ;
  input                                           std__pe45__lane28_strm0_data_valid  ;

  output                                          pe45__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane28_strm1_data_mask   ;
  input                                           std__pe45__lane28_strm1_data_valid  ;

  output                                          pe45__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane29_strm0_data_mask   ;
  input                                           std__pe45__lane29_strm0_data_valid  ;

  output                                          pe45__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane29_strm1_data_mask   ;
  input                                           std__pe45__lane29_strm1_data_valid  ;

  output                                          pe45__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane30_strm0_data_mask   ;
  input                                           std__pe45__lane30_strm0_data_valid  ;

  output                                          pe45__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane30_strm1_data_mask   ;
  input                                           std__pe45__lane30_strm1_data_valid  ;

  output                                          pe45__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane31_strm0_data_mask   ;
  input                                           std__pe45__lane31_strm0_data_valid  ;

  output                                          pe45__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe45__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe45__lane31_strm1_data_mask   ;
  input                                           std__pe45__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe46__peId                ;
  input                                         sys__pe46__allSynchronized     ;
  output                                        pe46__sys__thisSynchronized    ;
  output                                        pe46__sys__ready               ;
  output                                        pe46__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe46__oob_cntl            ;
  input                                         std__pe46__oob_valid           ;
  output                                        pe46__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe46__oob_type            ;
  output                                          pe46__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane0_strm0_data_mask   ;
  input                                           std__pe46__lane0_strm0_data_valid  ;

  output                                          pe46__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane0_strm1_data_mask   ;
  input                                           std__pe46__lane0_strm1_data_valid  ;

  output                                          pe46__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane1_strm0_data_mask   ;
  input                                           std__pe46__lane1_strm0_data_valid  ;

  output                                          pe46__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane1_strm1_data_mask   ;
  input                                           std__pe46__lane1_strm1_data_valid  ;

  output                                          pe46__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane2_strm0_data_mask   ;
  input                                           std__pe46__lane2_strm0_data_valid  ;

  output                                          pe46__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane2_strm1_data_mask   ;
  input                                           std__pe46__lane2_strm1_data_valid  ;

  output                                          pe46__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane3_strm0_data_mask   ;
  input                                           std__pe46__lane3_strm0_data_valid  ;

  output                                          pe46__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane3_strm1_data_mask   ;
  input                                           std__pe46__lane3_strm1_data_valid  ;

  output                                          pe46__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane4_strm0_data_mask   ;
  input                                           std__pe46__lane4_strm0_data_valid  ;

  output                                          pe46__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane4_strm1_data_mask   ;
  input                                           std__pe46__lane4_strm1_data_valid  ;

  output                                          pe46__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane5_strm0_data_mask   ;
  input                                           std__pe46__lane5_strm0_data_valid  ;

  output                                          pe46__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane5_strm1_data_mask   ;
  input                                           std__pe46__lane5_strm1_data_valid  ;

  output                                          pe46__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane6_strm0_data_mask   ;
  input                                           std__pe46__lane6_strm0_data_valid  ;

  output                                          pe46__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane6_strm1_data_mask   ;
  input                                           std__pe46__lane6_strm1_data_valid  ;

  output                                          pe46__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane7_strm0_data_mask   ;
  input                                           std__pe46__lane7_strm0_data_valid  ;

  output                                          pe46__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane7_strm1_data_mask   ;
  input                                           std__pe46__lane7_strm1_data_valid  ;

  output                                          pe46__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane8_strm0_data_mask   ;
  input                                           std__pe46__lane8_strm0_data_valid  ;

  output                                          pe46__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane8_strm1_data_mask   ;
  input                                           std__pe46__lane8_strm1_data_valid  ;

  output                                          pe46__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane9_strm0_data_mask   ;
  input                                           std__pe46__lane9_strm0_data_valid  ;

  output                                          pe46__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane9_strm1_data_mask   ;
  input                                           std__pe46__lane9_strm1_data_valid  ;

  output                                          pe46__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane10_strm0_data_mask   ;
  input                                           std__pe46__lane10_strm0_data_valid  ;

  output                                          pe46__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane10_strm1_data_mask   ;
  input                                           std__pe46__lane10_strm1_data_valid  ;

  output                                          pe46__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane11_strm0_data_mask   ;
  input                                           std__pe46__lane11_strm0_data_valid  ;

  output                                          pe46__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane11_strm1_data_mask   ;
  input                                           std__pe46__lane11_strm1_data_valid  ;

  output                                          pe46__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane12_strm0_data_mask   ;
  input                                           std__pe46__lane12_strm0_data_valid  ;

  output                                          pe46__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane12_strm1_data_mask   ;
  input                                           std__pe46__lane12_strm1_data_valid  ;

  output                                          pe46__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane13_strm0_data_mask   ;
  input                                           std__pe46__lane13_strm0_data_valid  ;

  output                                          pe46__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane13_strm1_data_mask   ;
  input                                           std__pe46__lane13_strm1_data_valid  ;

  output                                          pe46__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane14_strm0_data_mask   ;
  input                                           std__pe46__lane14_strm0_data_valid  ;

  output                                          pe46__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane14_strm1_data_mask   ;
  input                                           std__pe46__lane14_strm1_data_valid  ;

  output                                          pe46__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane15_strm0_data_mask   ;
  input                                           std__pe46__lane15_strm0_data_valid  ;

  output                                          pe46__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane15_strm1_data_mask   ;
  input                                           std__pe46__lane15_strm1_data_valid  ;

  output                                          pe46__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane16_strm0_data_mask   ;
  input                                           std__pe46__lane16_strm0_data_valid  ;

  output                                          pe46__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane16_strm1_data_mask   ;
  input                                           std__pe46__lane16_strm1_data_valid  ;

  output                                          pe46__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane17_strm0_data_mask   ;
  input                                           std__pe46__lane17_strm0_data_valid  ;

  output                                          pe46__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane17_strm1_data_mask   ;
  input                                           std__pe46__lane17_strm1_data_valid  ;

  output                                          pe46__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane18_strm0_data_mask   ;
  input                                           std__pe46__lane18_strm0_data_valid  ;

  output                                          pe46__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane18_strm1_data_mask   ;
  input                                           std__pe46__lane18_strm1_data_valid  ;

  output                                          pe46__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane19_strm0_data_mask   ;
  input                                           std__pe46__lane19_strm0_data_valid  ;

  output                                          pe46__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane19_strm1_data_mask   ;
  input                                           std__pe46__lane19_strm1_data_valid  ;

  output                                          pe46__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane20_strm0_data_mask   ;
  input                                           std__pe46__lane20_strm0_data_valid  ;

  output                                          pe46__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane20_strm1_data_mask   ;
  input                                           std__pe46__lane20_strm1_data_valid  ;

  output                                          pe46__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane21_strm0_data_mask   ;
  input                                           std__pe46__lane21_strm0_data_valid  ;

  output                                          pe46__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane21_strm1_data_mask   ;
  input                                           std__pe46__lane21_strm1_data_valid  ;

  output                                          pe46__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane22_strm0_data_mask   ;
  input                                           std__pe46__lane22_strm0_data_valid  ;

  output                                          pe46__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane22_strm1_data_mask   ;
  input                                           std__pe46__lane22_strm1_data_valid  ;

  output                                          pe46__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane23_strm0_data_mask   ;
  input                                           std__pe46__lane23_strm0_data_valid  ;

  output                                          pe46__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane23_strm1_data_mask   ;
  input                                           std__pe46__lane23_strm1_data_valid  ;

  output                                          pe46__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane24_strm0_data_mask   ;
  input                                           std__pe46__lane24_strm0_data_valid  ;

  output                                          pe46__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane24_strm1_data_mask   ;
  input                                           std__pe46__lane24_strm1_data_valid  ;

  output                                          pe46__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane25_strm0_data_mask   ;
  input                                           std__pe46__lane25_strm0_data_valid  ;

  output                                          pe46__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane25_strm1_data_mask   ;
  input                                           std__pe46__lane25_strm1_data_valid  ;

  output                                          pe46__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane26_strm0_data_mask   ;
  input                                           std__pe46__lane26_strm0_data_valid  ;

  output                                          pe46__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane26_strm1_data_mask   ;
  input                                           std__pe46__lane26_strm1_data_valid  ;

  output                                          pe46__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane27_strm0_data_mask   ;
  input                                           std__pe46__lane27_strm0_data_valid  ;

  output                                          pe46__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane27_strm1_data_mask   ;
  input                                           std__pe46__lane27_strm1_data_valid  ;

  output                                          pe46__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane28_strm0_data_mask   ;
  input                                           std__pe46__lane28_strm0_data_valid  ;

  output                                          pe46__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane28_strm1_data_mask   ;
  input                                           std__pe46__lane28_strm1_data_valid  ;

  output                                          pe46__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane29_strm0_data_mask   ;
  input                                           std__pe46__lane29_strm0_data_valid  ;

  output                                          pe46__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane29_strm1_data_mask   ;
  input                                           std__pe46__lane29_strm1_data_valid  ;

  output                                          pe46__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane30_strm0_data_mask   ;
  input                                           std__pe46__lane30_strm0_data_valid  ;

  output                                          pe46__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane30_strm1_data_mask   ;
  input                                           std__pe46__lane30_strm1_data_valid  ;

  output                                          pe46__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane31_strm0_data_mask   ;
  input                                           std__pe46__lane31_strm0_data_valid  ;

  output                                          pe46__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe46__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe46__lane31_strm1_data_mask   ;
  input                                           std__pe46__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe47__peId                ;
  input                                         sys__pe47__allSynchronized     ;
  output                                        pe47__sys__thisSynchronized    ;
  output                                        pe47__sys__ready               ;
  output                                        pe47__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe47__oob_cntl            ;
  input                                         std__pe47__oob_valid           ;
  output                                        pe47__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe47__oob_type            ;
  output                                          pe47__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane0_strm0_data_mask   ;
  input                                           std__pe47__lane0_strm0_data_valid  ;

  output                                          pe47__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane0_strm1_data_mask   ;
  input                                           std__pe47__lane0_strm1_data_valid  ;

  output                                          pe47__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane1_strm0_data_mask   ;
  input                                           std__pe47__lane1_strm0_data_valid  ;

  output                                          pe47__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane1_strm1_data_mask   ;
  input                                           std__pe47__lane1_strm1_data_valid  ;

  output                                          pe47__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane2_strm0_data_mask   ;
  input                                           std__pe47__lane2_strm0_data_valid  ;

  output                                          pe47__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane2_strm1_data_mask   ;
  input                                           std__pe47__lane2_strm1_data_valid  ;

  output                                          pe47__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane3_strm0_data_mask   ;
  input                                           std__pe47__lane3_strm0_data_valid  ;

  output                                          pe47__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane3_strm1_data_mask   ;
  input                                           std__pe47__lane3_strm1_data_valid  ;

  output                                          pe47__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane4_strm0_data_mask   ;
  input                                           std__pe47__lane4_strm0_data_valid  ;

  output                                          pe47__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane4_strm1_data_mask   ;
  input                                           std__pe47__lane4_strm1_data_valid  ;

  output                                          pe47__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane5_strm0_data_mask   ;
  input                                           std__pe47__lane5_strm0_data_valid  ;

  output                                          pe47__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane5_strm1_data_mask   ;
  input                                           std__pe47__lane5_strm1_data_valid  ;

  output                                          pe47__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane6_strm0_data_mask   ;
  input                                           std__pe47__lane6_strm0_data_valid  ;

  output                                          pe47__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane6_strm1_data_mask   ;
  input                                           std__pe47__lane6_strm1_data_valid  ;

  output                                          pe47__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane7_strm0_data_mask   ;
  input                                           std__pe47__lane7_strm0_data_valid  ;

  output                                          pe47__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane7_strm1_data_mask   ;
  input                                           std__pe47__lane7_strm1_data_valid  ;

  output                                          pe47__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane8_strm0_data_mask   ;
  input                                           std__pe47__lane8_strm0_data_valid  ;

  output                                          pe47__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane8_strm1_data_mask   ;
  input                                           std__pe47__lane8_strm1_data_valid  ;

  output                                          pe47__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane9_strm0_data_mask   ;
  input                                           std__pe47__lane9_strm0_data_valid  ;

  output                                          pe47__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane9_strm1_data_mask   ;
  input                                           std__pe47__lane9_strm1_data_valid  ;

  output                                          pe47__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane10_strm0_data_mask   ;
  input                                           std__pe47__lane10_strm0_data_valid  ;

  output                                          pe47__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane10_strm1_data_mask   ;
  input                                           std__pe47__lane10_strm1_data_valid  ;

  output                                          pe47__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane11_strm0_data_mask   ;
  input                                           std__pe47__lane11_strm0_data_valid  ;

  output                                          pe47__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane11_strm1_data_mask   ;
  input                                           std__pe47__lane11_strm1_data_valid  ;

  output                                          pe47__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane12_strm0_data_mask   ;
  input                                           std__pe47__lane12_strm0_data_valid  ;

  output                                          pe47__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane12_strm1_data_mask   ;
  input                                           std__pe47__lane12_strm1_data_valid  ;

  output                                          pe47__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane13_strm0_data_mask   ;
  input                                           std__pe47__lane13_strm0_data_valid  ;

  output                                          pe47__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane13_strm1_data_mask   ;
  input                                           std__pe47__lane13_strm1_data_valid  ;

  output                                          pe47__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane14_strm0_data_mask   ;
  input                                           std__pe47__lane14_strm0_data_valid  ;

  output                                          pe47__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane14_strm1_data_mask   ;
  input                                           std__pe47__lane14_strm1_data_valid  ;

  output                                          pe47__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane15_strm0_data_mask   ;
  input                                           std__pe47__lane15_strm0_data_valid  ;

  output                                          pe47__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane15_strm1_data_mask   ;
  input                                           std__pe47__lane15_strm1_data_valid  ;

  output                                          pe47__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane16_strm0_data_mask   ;
  input                                           std__pe47__lane16_strm0_data_valid  ;

  output                                          pe47__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane16_strm1_data_mask   ;
  input                                           std__pe47__lane16_strm1_data_valid  ;

  output                                          pe47__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane17_strm0_data_mask   ;
  input                                           std__pe47__lane17_strm0_data_valid  ;

  output                                          pe47__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane17_strm1_data_mask   ;
  input                                           std__pe47__lane17_strm1_data_valid  ;

  output                                          pe47__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane18_strm0_data_mask   ;
  input                                           std__pe47__lane18_strm0_data_valid  ;

  output                                          pe47__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane18_strm1_data_mask   ;
  input                                           std__pe47__lane18_strm1_data_valid  ;

  output                                          pe47__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane19_strm0_data_mask   ;
  input                                           std__pe47__lane19_strm0_data_valid  ;

  output                                          pe47__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane19_strm1_data_mask   ;
  input                                           std__pe47__lane19_strm1_data_valid  ;

  output                                          pe47__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane20_strm0_data_mask   ;
  input                                           std__pe47__lane20_strm0_data_valid  ;

  output                                          pe47__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane20_strm1_data_mask   ;
  input                                           std__pe47__lane20_strm1_data_valid  ;

  output                                          pe47__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane21_strm0_data_mask   ;
  input                                           std__pe47__lane21_strm0_data_valid  ;

  output                                          pe47__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane21_strm1_data_mask   ;
  input                                           std__pe47__lane21_strm1_data_valid  ;

  output                                          pe47__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane22_strm0_data_mask   ;
  input                                           std__pe47__lane22_strm0_data_valid  ;

  output                                          pe47__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane22_strm1_data_mask   ;
  input                                           std__pe47__lane22_strm1_data_valid  ;

  output                                          pe47__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane23_strm0_data_mask   ;
  input                                           std__pe47__lane23_strm0_data_valid  ;

  output                                          pe47__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane23_strm1_data_mask   ;
  input                                           std__pe47__lane23_strm1_data_valid  ;

  output                                          pe47__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane24_strm0_data_mask   ;
  input                                           std__pe47__lane24_strm0_data_valid  ;

  output                                          pe47__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane24_strm1_data_mask   ;
  input                                           std__pe47__lane24_strm1_data_valid  ;

  output                                          pe47__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane25_strm0_data_mask   ;
  input                                           std__pe47__lane25_strm0_data_valid  ;

  output                                          pe47__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane25_strm1_data_mask   ;
  input                                           std__pe47__lane25_strm1_data_valid  ;

  output                                          pe47__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane26_strm0_data_mask   ;
  input                                           std__pe47__lane26_strm0_data_valid  ;

  output                                          pe47__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane26_strm1_data_mask   ;
  input                                           std__pe47__lane26_strm1_data_valid  ;

  output                                          pe47__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane27_strm0_data_mask   ;
  input                                           std__pe47__lane27_strm0_data_valid  ;

  output                                          pe47__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane27_strm1_data_mask   ;
  input                                           std__pe47__lane27_strm1_data_valid  ;

  output                                          pe47__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane28_strm0_data_mask   ;
  input                                           std__pe47__lane28_strm0_data_valid  ;

  output                                          pe47__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane28_strm1_data_mask   ;
  input                                           std__pe47__lane28_strm1_data_valid  ;

  output                                          pe47__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane29_strm0_data_mask   ;
  input                                           std__pe47__lane29_strm0_data_valid  ;

  output                                          pe47__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane29_strm1_data_mask   ;
  input                                           std__pe47__lane29_strm1_data_valid  ;

  output                                          pe47__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane30_strm0_data_mask   ;
  input                                           std__pe47__lane30_strm0_data_valid  ;

  output                                          pe47__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane30_strm1_data_mask   ;
  input                                           std__pe47__lane30_strm1_data_valid  ;

  output                                          pe47__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane31_strm0_data_mask   ;
  input                                           std__pe47__lane31_strm0_data_valid  ;

  output                                          pe47__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe47__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe47__lane31_strm1_data_mask   ;
  input                                           std__pe47__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe48__peId                ;
  input                                         sys__pe48__allSynchronized     ;
  output                                        pe48__sys__thisSynchronized    ;
  output                                        pe48__sys__ready               ;
  output                                        pe48__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe48__oob_cntl            ;
  input                                         std__pe48__oob_valid           ;
  output                                        pe48__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe48__oob_type            ;
  output                                          pe48__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane0_strm0_data_mask   ;
  input                                           std__pe48__lane0_strm0_data_valid  ;

  output                                          pe48__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane0_strm1_data_mask   ;
  input                                           std__pe48__lane0_strm1_data_valid  ;

  output                                          pe48__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane1_strm0_data_mask   ;
  input                                           std__pe48__lane1_strm0_data_valid  ;

  output                                          pe48__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane1_strm1_data_mask   ;
  input                                           std__pe48__lane1_strm1_data_valid  ;

  output                                          pe48__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane2_strm0_data_mask   ;
  input                                           std__pe48__lane2_strm0_data_valid  ;

  output                                          pe48__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane2_strm1_data_mask   ;
  input                                           std__pe48__lane2_strm1_data_valid  ;

  output                                          pe48__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane3_strm0_data_mask   ;
  input                                           std__pe48__lane3_strm0_data_valid  ;

  output                                          pe48__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane3_strm1_data_mask   ;
  input                                           std__pe48__lane3_strm1_data_valid  ;

  output                                          pe48__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane4_strm0_data_mask   ;
  input                                           std__pe48__lane4_strm0_data_valid  ;

  output                                          pe48__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane4_strm1_data_mask   ;
  input                                           std__pe48__lane4_strm1_data_valid  ;

  output                                          pe48__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane5_strm0_data_mask   ;
  input                                           std__pe48__lane5_strm0_data_valid  ;

  output                                          pe48__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane5_strm1_data_mask   ;
  input                                           std__pe48__lane5_strm1_data_valid  ;

  output                                          pe48__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane6_strm0_data_mask   ;
  input                                           std__pe48__lane6_strm0_data_valid  ;

  output                                          pe48__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane6_strm1_data_mask   ;
  input                                           std__pe48__lane6_strm1_data_valid  ;

  output                                          pe48__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane7_strm0_data_mask   ;
  input                                           std__pe48__lane7_strm0_data_valid  ;

  output                                          pe48__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane7_strm1_data_mask   ;
  input                                           std__pe48__lane7_strm1_data_valid  ;

  output                                          pe48__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane8_strm0_data_mask   ;
  input                                           std__pe48__lane8_strm0_data_valid  ;

  output                                          pe48__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane8_strm1_data_mask   ;
  input                                           std__pe48__lane8_strm1_data_valid  ;

  output                                          pe48__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane9_strm0_data_mask   ;
  input                                           std__pe48__lane9_strm0_data_valid  ;

  output                                          pe48__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane9_strm1_data_mask   ;
  input                                           std__pe48__lane9_strm1_data_valid  ;

  output                                          pe48__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane10_strm0_data_mask   ;
  input                                           std__pe48__lane10_strm0_data_valid  ;

  output                                          pe48__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane10_strm1_data_mask   ;
  input                                           std__pe48__lane10_strm1_data_valid  ;

  output                                          pe48__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane11_strm0_data_mask   ;
  input                                           std__pe48__lane11_strm0_data_valid  ;

  output                                          pe48__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane11_strm1_data_mask   ;
  input                                           std__pe48__lane11_strm1_data_valid  ;

  output                                          pe48__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane12_strm0_data_mask   ;
  input                                           std__pe48__lane12_strm0_data_valid  ;

  output                                          pe48__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane12_strm1_data_mask   ;
  input                                           std__pe48__lane12_strm1_data_valid  ;

  output                                          pe48__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane13_strm0_data_mask   ;
  input                                           std__pe48__lane13_strm0_data_valid  ;

  output                                          pe48__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane13_strm1_data_mask   ;
  input                                           std__pe48__lane13_strm1_data_valid  ;

  output                                          pe48__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane14_strm0_data_mask   ;
  input                                           std__pe48__lane14_strm0_data_valid  ;

  output                                          pe48__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane14_strm1_data_mask   ;
  input                                           std__pe48__lane14_strm1_data_valid  ;

  output                                          pe48__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane15_strm0_data_mask   ;
  input                                           std__pe48__lane15_strm0_data_valid  ;

  output                                          pe48__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane15_strm1_data_mask   ;
  input                                           std__pe48__lane15_strm1_data_valid  ;

  output                                          pe48__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane16_strm0_data_mask   ;
  input                                           std__pe48__lane16_strm0_data_valid  ;

  output                                          pe48__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane16_strm1_data_mask   ;
  input                                           std__pe48__lane16_strm1_data_valid  ;

  output                                          pe48__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane17_strm0_data_mask   ;
  input                                           std__pe48__lane17_strm0_data_valid  ;

  output                                          pe48__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane17_strm1_data_mask   ;
  input                                           std__pe48__lane17_strm1_data_valid  ;

  output                                          pe48__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane18_strm0_data_mask   ;
  input                                           std__pe48__lane18_strm0_data_valid  ;

  output                                          pe48__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane18_strm1_data_mask   ;
  input                                           std__pe48__lane18_strm1_data_valid  ;

  output                                          pe48__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane19_strm0_data_mask   ;
  input                                           std__pe48__lane19_strm0_data_valid  ;

  output                                          pe48__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane19_strm1_data_mask   ;
  input                                           std__pe48__lane19_strm1_data_valid  ;

  output                                          pe48__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane20_strm0_data_mask   ;
  input                                           std__pe48__lane20_strm0_data_valid  ;

  output                                          pe48__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane20_strm1_data_mask   ;
  input                                           std__pe48__lane20_strm1_data_valid  ;

  output                                          pe48__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane21_strm0_data_mask   ;
  input                                           std__pe48__lane21_strm0_data_valid  ;

  output                                          pe48__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane21_strm1_data_mask   ;
  input                                           std__pe48__lane21_strm1_data_valid  ;

  output                                          pe48__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane22_strm0_data_mask   ;
  input                                           std__pe48__lane22_strm0_data_valid  ;

  output                                          pe48__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane22_strm1_data_mask   ;
  input                                           std__pe48__lane22_strm1_data_valid  ;

  output                                          pe48__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane23_strm0_data_mask   ;
  input                                           std__pe48__lane23_strm0_data_valid  ;

  output                                          pe48__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane23_strm1_data_mask   ;
  input                                           std__pe48__lane23_strm1_data_valid  ;

  output                                          pe48__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane24_strm0_data_mask   ;
  input                                           std__pe48__lane24_strm0_data_valid  ;

  output                                          pe48__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane24_strm1_data_mask   ;
  input                                           std__pe48__lane24_strm1_data_valid  ;

  output                                          pe48__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane25_strm0_data_mask   ;
  input                                           std__pe48__lane25_strm0_data_valid  ;

  output                                          pe48__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane25_strm1_data_mask   ;
  input                                           std__pe48__lane25_strm1_data_valid  ;

  output                                          pe48__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane26_strm0_data_mask   ;
  input                                           std__pe48__lane26_strm0_data_valid  ;

  output                                          pe48__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane26_strm1_data_mask   ;
  input                                           std__pe48__lane26_strm1_data_valid  ;

  output                                          pe48__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane27_strm0_data_mask   ;
  input                                           std__pe48__lane27_strm0_data_valid  ;

  output                                          pe48__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane27_strm1_data_mask   ;
  input                                           std__pe48__lane27_strm1_data_valid  ;

  output                                          pe48__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane28_strm0_data_mask   ;
  input                                           std__pe48__lane28_strm0_data_valid  ;

  output                                          pe48__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane28_strm1_data_mask   ;
  input                                           std__pe48__lane28_strm1_data_valid  ;

  output                                          pe48__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane29_strm0_data_mask   ;
  input                                           std__pe48__lane29_strm0_data_valid  ;

  output                                          pe48__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane29_strm1_data_mask   ;
  input                                           std__pe48__lane29_strm1_data_valid  ;

  output                                          pe48__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane30_strm0_data_mask   ;
  input                                           std__pe48__lane30_strm0_data_valid  ;

  output                                          pe48__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane30_strm1_data_mask   ;
  input                                           std__pe48__lane30_strm1_data_valid  ;

  output                                          pe48__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane31_strm0_data_mask   ;
  input                                           std__pe48__lane31_strm0_data_valid  ;

  output                                          pe48__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe48__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe48__lane31_strm1_data_mask   ;
  input                                           std__pe48__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe49__peId                ;
  input                                         sys__pe49__allSynchronized     ;
  output                                        pe49__sys__thisSynchronized    ;
  output                                        pe49__sys__ready               ;
  output                                        pe49__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe49__oob_cntl            ;
  input                                         std__pe49__oob_valid           ;
  output                                        pe49__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe49__oob_type            ;
  output                                          pe49__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane0_strm0_data_mask   ;
  input                                           std__pe49__lane0_strm0_data_valid  ;

  output                                          pe49__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane0_strm1_data_mask   ;
  input                                           std__pe49__lane0_strm1_data_valid  ;

  output                                          pe49__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane1_strm0_data_mask   ;
  input                                           std__pe49__lane1_strm0_data_valid  ;

  output                                          pe49__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane1_strm1_data_mask   ;
  input                                           std__pe49__lane1_strm1_data_valid  ;

  output                                          pe49__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane2_strm0_data_mask   ;
  input                                           std__pe49__lane2_strm0_data_valid  ;

  output                                          pe49__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane2_strm1_data_mask   ;
  input                                           std__pe49__lane2_strm1_data_valid  ;

  output                                          pe49__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane3_strm0_data_mask   ;
  input                                           std__pe49__lane3_strm0_data_valid  ;

  output                                          pe49__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane3_strm1_data_mask   ;
  input                                           std__pe49__lane3_strm1_data_valid  ;

  output                                          pe49__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane4_strm0_data_mask   ;
  input                                           std__pe49__lane4_strm0_data_valid  ;

  output                                          pe49__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane4_strm1_data_mask   ;
  input                                           std__pe49__lane4_strm1_data_valid  ;

  output                                          pe49__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane5_strm0_data_mask   ;
  input                                           std__pe49__lane5_strm0_data_valid  ;

  output                                          pe49__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane5_strm1_data_mask   ;
  input                                           std__pe49__lane5_strm1_data_valid  ;

  output                                          pe49__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane6_strm0_data_mask   ;
  input                                           std__pe49__lane6_strm0_data_valid  ;

  output                                          pe49__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane6_strm1_data_mask   ;
  input                                           std__pe49__lane6_strm1_data_valid  ;

  output                                          pe49__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane7_strm0_data_mask   ;
  input                                           std__pe49__lane7_strm0_data_valid  ;

  output                                          pe49__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane7_strm1_data_mask   ;
  input                                           std__pe49__lane7_strm1_data_valid  ;

  output                                          pe49__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane8_strm0_data_mask   ;
  input                                           std__pe49__lane8_strm0_data_valid  ;

  output                                          pe49__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane8_strm1_data_mask   ;
  input                                           std__pe49__lane8_strm1_data_valid  ;

  output                                          pe49__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane9_strm0_data_mask   ;
  input                                           std__pe49__lane9_strm0_data_valid  ;

  output                                          pe49__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane9_strm1_data_mask   ;
  input                                           std__pe49__lane9_strm1_data_valid  ;

  output                                          pe49__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane10_strm0_data_mask   ;
  input                                           std__pe49__lane10_strm0_data_valid  ;

  output                                          pe49__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane10_strm1_data_mask   ;
  input                                           std__pe49__lane10_strm1_data_valid  ;

  output                                          pe49__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane11_strm0_data_mask   ;
  input                                           std__pe49__lane11_strm0_data_valid  ;

  output                                          pe49__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane11_strm1_data_mask   ;
  input                                           std__pe49__lane11_strm1_data_valid  ;

  output                                          pe49__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane12_strm0_data_mask   ;
  input                                           std__pe49__lane12_strm0_data_valid  ;

  output                                          pe49__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane12_strm1_data_mask   ;
  input                                           std__pe49__lane12_strm1_data_valid  ;

  output                                          pe49__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane13_strm0_data_mask   ;
  input                                           std__pe49__lane13_strm0_data_valid  ;

  output                                          pe49__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane13_strm1_data_mask   ;
  input                                           std__pe49__lane13_strm1_data_valid  ;

  output                                          pe49__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane14_strm0_data_mask   ;
  input                                           std__pe49__lane14_strm0_data_valid  ;

  output                                          pe49__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane14_strm1_data_mask   ;
  input                                           std__pe49__lane14_strm1_data_valid  ;

  output                                          pe49__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane15_strm0_data_mask   ;
  input                                           std__pe49__lane15_strm0_data_valid  ;

  output                                          pe49__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane15_strm1_data_mask   ;
  input                                           std__pe49__lane15_strm1_data_valid  ;

  output                                          pe49__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane16_strm0_data_mask   ;
  input                                           std__pe49__lane16_strm0_data_valid  ;

  output                                          pe49__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane16_strm1_data_mask   ;
  input                                           std__pe49__lane16_strm1_data_valid  ;

  output                                          pe49__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane17_strm0_data_mask   ;
  input                                           std__pe49__lane17_strm0_data_valid  ;

  output                                          pe49__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane17_strm1_data_mask   ;
  input                                           std__pe49__lane17_strm1_data_valid  ;

  output                                          pe49__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane18_strm0_data_mask   ;
  input                                           std__pe49__lane18_strm0_data_valid  ;

  output                                          pe49__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane18_strm1_data_mask   ;
  input                                           std__pe49__lane18_strm1_data_valid  ;

  output                                          pe49__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane19_strm0_data_mask   ;
  input                                           std__pe49__lane19_strm0_data_valid  ;

  output                                          pe49__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane19_strm1_data_mask   ;
  input                                           std__pe49__lane19_strm1_data_valid  ;

  output                                          pe49__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane20_strm0_data_mask   ;
  input                                           std__pe49__lane20_strm0_data_valid  ;

  output                                          pe49__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane20_strm1_data_mask   ;
  input                                           std__pe49__lane20_strm1_data_valid  ;

  output                                          pe49__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane21_strm0_data_mask   ;
  input                                           std__pe49__lane21_strm0_data_valid  ;

  output                                          pe49__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane21_strm1_data_mask   ;
  input                                           std__pe49__lane21_strm1_data_valid  ;

  output                                          pe49__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane22_strm0_data_mask   ;
  input                                           std__pe49__lane22_strm0_data_valid  ;

  output                                          pe49__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane22_strm1_data_mask   ;
  input                                           std__pe49__lane22_strm1_data_valid  ;

  output                                          pe49__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane23_strm0_data_mask   ;
  input                                           std__pe49__lane23_strm0_data_valid  ;

  output                                          pe49__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane23_strm1_data_mask   ;
  input                                           std__pe49__lane23_strm1_data_valid  ;

  output                                          pe49__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane24_strm0_data_mask   ;
  input                                           std__pe49__lane24_strm0_data_valid  ;

  output                                          pe49__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane24_strm1_data_mask   ;
  input                                           std__pe49__lane24_strm1_data_valid  ;

  output                                          pe49__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane25_strm0_data_mask   ;
  input                                           std__pe49__lane25_strm0_data_valid  ;

  output                                          pe49__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane25_strm1_data_mask   ;
  input                                           std__pe49__lane25_strm1_data_valid  ;

  output                                          pe49__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane26_strm0_data_mask   ;
  input                                           std__pe49__lane26_strm0_data_valid  ;

  output                                          pe49__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane26_strm1_data_mask   ;
  input                                           std__pe49__lane26_strm1_data_valid  ;

  output                                          pe49__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane27_strm0_data_mask   ;
  input                                           std__pe49__lane27_strm0_data_valid  ;

  output                                          pe49__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane27_strm1_data_mask   ;
  input                                           std__pe49__lane27_strm1_data_valid  ;

  output                                          pe49__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane28_strm0_data_mask   ;
  input                                           std__pe49__lane28_strm0_data_valid  ;

  output                                          pe49__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane28_strm1_data_mask   ;
  input                                           std__pe49__lane28_strm1_data_valid  ;

  output                                          pe49__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane29_strm0_data_mask   ;
  input                                           std__pe49__lane29_strm0_data_valid  ;

  output                                          pe49__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane29_strm1_data_mask   ;
  input                                           std__pe49__lane29_strm1_data_valid  ;

  output                                          pe49__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane30_strm0_data_mask   ;
  input                                           std__pe49__lane30_strm0_data_valid  ;

  output                                          pe49__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane30_strm1_data_mask   ;
  input                                           std__pe49__lane30_strm1_data_valid  ;

  output                                          pe49__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane31_strm0_data_mask   ;
  input                                           std__pe49__lane31_strm0_data_valid  ;

  output                                          pe49__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe49__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe49__lane31_strm1_data_mask   ;
  input                                           std__pe49__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe50__peId                ;
  input                                         sys__pe50__allSynchronized     ;
  output                                        pe50__sys__thisSynchronized    ;
  output                                        pe50__sys__ready               ;
  output                                        pe50__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe50__oob_cntl            ;
  input                                         std__pe50__oob_valid           ;
  output                                        pe50__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe50__oob_type            ;
  output                                          pe50__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane0_strm0_data_mask   ;
  input                                           std__pe50__lane0_strm0_data_valid  ;

  output                                          pe50__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane0_strm1_data_mask   ;
  input                                           std__pe50__lane0_strm1_data_valid  ;

  output                                          pe50__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane1_strm0_data_mask   ;
  input                                           std__pe50__lane1_strm0_data_valid  ;

  output                                          pe50__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane1_strm1_data_mask   ;
  input                                           std__pe50__lane1_strm1_data_valid  ;

  output                                          pe50__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane2_strm0_data_mask   ;
  input                                           std__pe50__lane2_strm0_data_valid  ;

  output                                          pe50__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane2_strm1_data_mask   ;
  input                                           std__pe50__lane2_strm1_data_valid  ;

  output                                          pe50__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane3_strm0_data_mask   ;
  input                                           std__pe50__lane3_strm0_data_valid  ;

  output                                          pe50__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane3_strm1_data_mask   ;
  input                                           std__pe50__lane3_strm1_data_valid  ;

  output                                          pe50__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane4_strm0_data_mask   ;
  input                                           std__pe50__lane4_strm0_data_valid  ;

  output                                          pe50__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane4_strm1_data_mask   ;
  input                                           std__pe50__lane4_strm1_data_valid  ;

  output                                          pe50__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane5_strm0_data_mask   ;
  input                                           std__pe50__lane5_strm0_data_valid  ;

  output                                          pe50__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane5_strm1_data_mask   ;
  input                                           std__pe50__lane5_strm1_data_valid  ;

  output                                          pe50__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane6_strm0_data_mask   ;
  input                                           std__pe50__lane6_strm0_data_valid  ;

  output                                          pe50__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane6_strm1_data_mask   ;
  input                                           std__pe50__lane6_strm1_data_valid  ;

  output                                          pe50__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane7_strm0_data_mask   ;
  input                                           std__pe50__lane7_strm0_data_valid  ;

  output                                          pe50__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane7_strm1_data_mask   ;
  input                                           std__pe50__lane7_strm1_data_valid  ;

  output                                          pe50__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane8_strm0_data_mask   ;
  input                                           std__pe50__lane8_strm0_data_valid  ;

  output                                          pe50__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane8_strm1_data_mask   ;
  input                                           std__pe50__lane8_strm1_data_valid  ;

  output                                          pe50__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane9_strm0_data_mask   ;
  input                                           std__pe50__lane9_strm0_data_valid  ;

  output                                          pe50__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane9_strm1_data_mask   ;
  input                                           std__pe50__lane9_strm1_data_valid  ;

  output                                          pe50__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane10_strm0_data_mask   ;
  input                                           std__pe50__lane10_strm0_data_valid  ;

  output                                          pe50__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane10_strm1_data_mask   ;
  input                                           std__pe50__lane10_strm1_data_valid  ;

  output                                          pe50__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane11_strm0_data_mask   ;
  input                                           std__pe50__lane11_strm0_data_valid  ;

  output                                          pe50__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane11_strm1_data_mask   ;
  input                                           std__pe50__lane11_strm1_data_valid  ;

  output                                          pe50__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane12_strm0_data_mask   ;
  input                                           std__pe50__lane12_strm0_data_valid  ;

  output                                          pe50__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane12_strm1_data_mask   ;
  input                                           std__pe50__lane12_strm1_data_valid  ;

  output                                          pe50__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane13_strm0_data_mask   ;
  input                                           std__pe50__lane13_strm0_data_valid  ;

  output                                          pe50__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane13_strm1_data_mask   ;
  input                                           std__pe50__lane13_strm1_data_valid  ;

  output                                          pe50__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane14_strm0_data_mask   ;
  input                                           std__pe50__lane14_strm0_data_valid  ;

  output                                          pe50__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane14_strm1_data_mask   ;
  input                                           std__pe50__lane14_strm1_data_valid  ;

  output                                          pe50__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane15_strm0_data_mask   ;
  input                                           std__pe50__lane15_strm0_data_valid  ;

  output                                          pe50__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane15_strm1_data_mask   ;
  input                                           std__pe50__lane15_strm1_data_valid  ;

  output                                          pe50__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane16_strm0_data_mask   ;
  input                                           std__pe50__lane16_strm0_data_valid  ;

  output                                          pe50__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane16_strm1_data_mask   ;
  input                                           std__pe50__lane16_strm1_data_valid  ;

  output                                          pe50__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane17_strm0_data_mask   ;
  input                                           std__pe50__lane17_strm0_data_valid  ;

  output                                          pe50__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane17_strm1_data_mask   ;
  input                                           std__pe50__lane17_strm1_data_valid  ;

  output                                          pe50__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane18_strm0_data_mask   ;
  input                                           std__pe50__lane18_strm0_data_valid  ;

  output                                          pe50__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane18_strm1_data_mask   ;
  input                                           std__pe50__lane18_strm1_data_valid  ;

  output                                          pe50__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane19_strm0_data_mask   ;
  input                                           std__pe50__lane19_strm0_data_valid  ;

  output                                          pe50__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane19_strm1_data_mask   ;
  input                                           std__pe50__lane19_strm1_data_valid  ;

  output                                          pe50__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane20_strm0_data_mask   ;
  input                                           std__pe50__lane20_strm0_data_valid  ;

  output                                          pe50__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane20_strm1_data_mask   ;
  input                                           std__pe50__lane20_strm1_data_valid  ;

  output                                          pe50__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane21_strm0_data_mask   ;
  input                                           std__pe50__lane21_strm0_data_valid  ;

  output                                          pe50__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane21_strm1_data_mask   ;
  input                                           std__pe50__lane21_strm1_data_valid  ;

  output                                          pe50__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane22_strm0_data_mask   ;
  input                                           std__pe50__lane22_strm0_data_valid  ;

  output                                          pe50__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane22_strm1_data_mask   ;
  input                                           std__pe50__lane22_strm1_data_valid  ;

  output                                          pe50__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane23_strm0_data_mask   ;
  input                                           std__pe50__lane23_strm0_data_valid  ;

  output                                          pe50__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane23_strm1_data_mask   ;
  input                                           std__pe50__lane23_strm1_data_valid  ;

  output                                          pe50__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane24_strm0_data_mask   ;
  input                                           std__pe50__lane24_strm0_data_valid  ;

  output                                          pe50__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane24_strm1_data_mask   ;
  input                                           std__pe50__lane24_strm1_data_valid  ;

  output                                          pe50__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane25_strm0_data_mask   ;
  input                                           std__pe50__lane25_strm0_data_valid  ;

  output                                          pe50__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane25_strm1_data_mask   ;
  input                                           std__pe50__lane25_strm1_data_valid  ;

  output                                          pe50__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane26_strm0_data_mask   ;
  input                                           std__pe50__lane26_strm0_data_valid  ;

  output                                          pe50__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane26_strm1_data_mask   ;
  input                                           std__pe50__lane26_strm1_data_valid  ;

  output                                          pe50__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane27_strm0_data_mask   ;
  input                                           std__pe50__lane27_strm0_data_valid  ;

  output                                          pe50__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane27_strm1_data_mask   ;
  input                                           std__pe50__lane27_strm1_data_valid  ;

  output                                          pe50__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane28_strm0_data_mask   ;
  input                                           std__pe50__lane28_strm0_data_valid  ;

  output                                          pe50__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane28_strm1_data_mask   ;
  input                                           std__pe50__lane28_strm1_data_valid  ;

  output                                          pe50__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane29_strm0_data_mask   ;
  input                                           std__pe50__lane29_strm0_data_valid  ;

  output                                          pe50__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane29_strm1_data_mask   ;
  input                                           std__pe50__lane29_strm1_data_valid  ;

  output                                          pe50__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane30_strm0_data_mask   ;
  input                                           std__pe50__lane30_strm0_data_valid  ;

  output                                          pe50__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane30_strm1_data_mask   ;
  input                                           std__pe50__lane30_strm1_data_valid  ;

  output                                          pe50__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane31_strm0_data_mask   ;
  input                                           std__pe50__lane31_strm0_data_valid  ;

  output                                          pe50__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe50__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe50__lane31_strm1_data_mask   ;
  input                                           std__pe50__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe51__peId                ;
  input                                         sys__pe51__allSynchronized     ;
  output                                        pe51__sys__thisSynchronized    ;
  output                                        pe51__sys__ready               ;
  output                                        pe51__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe51__oob_cntl            ;
  input                                         std__pe51__oob_valid           ;
  output                                        pe51__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe51__oob_type            ;
  output                                          pe51__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane0_strm0_data_mask   ;
  input                                           std__pe51__lane0_strm0_data_valid  ;

  output                                          pe51__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane0_strm1_data_mask   ;
  input                                           std__pe51__lane0_strm1_data_valid  ;

  output                                          pe51__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane1_strm0_data_mask   ;
  input                                           std__pe51__lane1_strm0_data_valid  ;

  output                                          pe51__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane1_strm1_data_mask   ;
  input                                           std__pe51__lane1_strm1_data_valid  ;

  output                                          pe51__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane2_strm0_data_mask   ;
  input                                           std__pe51__lane2_strm0_data_valid  ;

  output                                          pe51__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane2_strm1_data_mask   ;
  input                                           std__pe51__lane2_strm1_data_valid  ;

  output                                          pe51__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane3_strm0_data_mask   ;
  input                                           std__pe51__lane3_strm0_data_valid  ;

  output                                          pe51__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane3_strm1_data_mask   ;
  input                                           std__pe51__lane3_strm1_data_valid  ;

  output                                          pe51__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane4_strm0_data_mask   ;
  input                                           std__pe51__lane4_strm0_data_valid  ;

  output                                          pe51__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane4_strm1_data_mask   ;
  input                                           std__pe51__lane4_strm1_data_valid  ;

  output                                          pe51__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane5_strm0_data_mask   ;
  input                                           std__pe51__lane5_strm0_data_valid  ;

  output                                          pe51__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane5_strm1_data_mask   ;
  input                                           std__pe51__lane5_strm1_data_valid  ;

  output                                          pe51__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane6_strm0_data_mask   ;
  input                                           std__pe51__lane6_strm0_data_valid  ;

  output                                          pe51__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane6_strm1_data_mask   ;
  input                                           std__pe51__lane6_strm1_data_valid  ;

  output                                          pe51__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane7_strm0_data_mask   ;
  input                                           std__pe51__lane7_strm0_data_valid  ;

  output                                          pe51__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane7_strm1_data_mask   ;
  input                                           std__pe51__lane7_strm1_data_valid  ;

  output                                          pe51__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane8_strm0_data_mask   ;
  input                                           std__pe51__lane8_strm0_data_valid  ;

  output                                          pe51__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane8_strm1_data_mask   ;
  input                                           std__pe51__lane8_strm1_data_valid  ;

  output                                          pe51__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane9_strm0_data_mask   ;
  input                                           std__pe51__lane9_strm0_data_valid  ;

  output                                          pe51__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane9_strm1_data_mask   ;
  input                                           std__pe51__lane9_strm1_data_valid  ;

  output                                          pe51__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane10_strm0_data_mask   ;
  input                                           std__pe51__lane10_strm0_data_valid  ;

  output                                          pe51__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane10_strm1_data_mask   ;
  input                                           std__pe51__lane10_strm1_data_valid  ;

  output                                          pe51__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane11_strm0_data_mask   ;
  input                                           std__pe51__lane11_strm0_data_valid  ;

  output                                          pe51__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane11_strm1_data_mask   ;
  input                                           std__pe51__lane11_strm1_data_valid  ;

  output                                          pe51__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane12_strm0_data_mask   ;
  input                                           std__pe51__lane12_strm0_data_valid  ;

  output                                          pe51__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane12_strm1_data_mask   ;
  input                                           std__pe51__lane12_strm1_data_valid  ;

  output                                          pe51__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane13_strm0_data_mask   ;
  input                                           std__pe51__lane13_strm0_data_valid  ;

  output                                          pe51__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane13_strm1_data_mask   ;
  input                                           std__pe51__lane13_strm1_data_valid  ;

  output                                          pe51__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane14_strm0_data_mask   ;
  input                                           std__pe51__lane14_strm0_data_valid  ;

  output                                          pe51__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane14_strm1_data_mask   ;
  input                                           std__pe51__lane14_strm1_data_valid  ;

  output                                          pe51__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane15_strm0_data_mask   ;
  input                                           std__pe51__lane15_strm0_data_valid  ;

  output                                          pe51__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane15_strm1_data_mask   ;
  input                                           std__pe51__lane15_strm1_data_valid  ;

  output                                          pe51__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane16_strm0_data_mask   ;
  input                                           std__pe51__lane16_strm0_data_valid  ;

  output                                          pe51__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane16_strm1_data_mask   ;
  input                                           std__pe51__lane16_strm1_data_valid  ;

  output                                          pe51__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane17_strm0_data_mask   ;
  input                                           std__pe51__lane17_strm0_data_valid  ;

  output                                          pe51__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane17_strm1_data_mask   ;
  input                                           std__pe51__lane17_strm1_data_valid  ;

  output                                          pe51__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane18_strm0_data_mask   ;
  input                                           std__pe51__lane18_strm0_data_valid  ;

  output                                          pe51__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane18_strm1_data_mask   ;
  input                                           std__pe51__lane18_strm1_data_valid  ;

  output                                          pe51__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane19_strm0_data_mask   ;
  input                                           std__pe51__lane19_strm0_data_valid  ;

  output                                          pe51__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane19_strm1_data_mask   ;
  input                                           std__pe51__lane19_strm1_data_valid  ;

  output                                          pe51__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane20_strm0_data_mask   ;
  input                                           std__pe51__lane20_strm0_data_valid  ;

  output                                          pe51__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane20_strm1_data_mask   ;
  input                                           std__pe51__lane20_strm1_data_valid  ;

  output                                          pe51__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane21_strm0_data_mask   ;
  input                                           std__pe51__lane21_strm0_data_valid  ;

  output                                          pe51__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane21_strm1_data_mask   ;
  input                                           std__pe51__lane21_strm1_data_valid  ;

  output                                          pe51__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane22_strm0_data_mask   ;
  input                                           std__pe51__lane22_strm0_data_valid  ;

  output                                          pe51__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane22_strm1_data_mask   ;
  input                                           std__pe51__lane22_strm1_data_valid  ;

  output                                          pe51__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane23_strm0_data_mask   ;
  input                                           std__pe51__lane23_strm0_data_valid  ;

  output                                          pe51__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane23_strm1_data_mask   ;
  input                                           std__pe51__lane23_strm1_data_valid  ;

  output                                          pe51__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane24_strm0_data_mask   ;
  input                                           std__pe51__lane24_strm0_data_valid  ;

  output                                          pe51__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane24_strm1_data_mask   ;
  input                                           std__pe51__lane24_strm1_data_valid  ;

  output                                          pe51__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane25_strm0_data_mask   ;
  input                                           std__pe51__lane25_strm0_data_valid  ;

  output                                          pe51__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane25_strm1_data_mask   ;
  input                                           std__pe51__lane25_strm1_data_valid  ;

  output                                          pe51__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane26_strm0_data_mask   ;
  input                                           std__pe51__lane26_strm0_data_valid  ;

  output                                          pe51__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane26_strm1_data_mask   ;
  input                                           std__pe51__lane26_strm1_data_valid  ;

  output                                          pe51__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane27_strm0_data_mask   ;
  input                                           std__pe51__lane27_strm0_data_valid  ;

  output                                          pe51__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane27_strm1_data_mask   ;
  input                                           std__pe51__lane27_strm1_data_valid  ;

  output                                          pe51__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane28_strm0_data_mask   ;
  input                                           std__pe51__lane28_strm0_data_valid  ;

  output                                          pe51__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane28_strm1_data_mask   ;
  input                                           std__pe51__lane28_strm1_data_valid  ;

  output                                          pe51__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane29_strm0_data_mask   ;
  input                                           std__pe51__lane29_strm0_data_valid  ;

  output                                          pe51__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane29_strm1_data_mask   ;
  input                                           std__pe51__lane29_strm1_data_valid  ;

  output                                          pe51__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane30_strm0_data_mask   ;
  input                                           std__pe51__lane30_strm0_data_valid  ;

  output                                          pe51__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane30_strm1_data_mask   ;
  input                                           std__pe51__lane30_strm1_data_valid  ;

  output                                          pe51__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane31_strm0_data_mask   ;
  input                                           std__pe51__lane31_strm0_data_valid  ;

  output                                          pe51__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe51__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe51__lane31_strm1_data_mask   ;
  input                                           std__pe51__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe52__peId                ;
  input                                         sys__pe52__allSynchronized     ;
  output                                        pe52__sys__thisSynchronized    ;
  output                                        pe52__sys__ready               ;
  output                                        pe52__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe52__oob_cntl            ;
  input                                         std__pe52__oob_valid           ;
  output                                        pe52__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe52__oob_type            ;
  output                                          pe52__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane0_strm0_data_mask   ;
  input                                           std__pe52__lane0_strm0_data_valid  ;

  output                                          pe52__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane0_strm1_data_mask   ;
  input                                           std__pe52__lane0_strm1_data_valid  ;

  output                                          pe52__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane1_strm0_data_mask   ;
  input                                           std__pe52__lane1_strm0_data_valid  ;

  output                                          pe52__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane1_strm1_data_mask   ;
  input                                           std__pe52__lane1_strm1_data_valid  ;

  output                                          pe52__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane2_strm0_data_mask   ;
  input                                           std__pe52__lane2_strm0_data_valid  ;

  output                                          pe52__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane2_strm1_data_mask   ;
  input                                           std__pe52__lane2_strm1_data_valid  ;

  output                                          pe52__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane3_strm0_data_mask   ;
  input                                           std__pe52__lane3_strm0_data_valid  ;

  output                                          pe52__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane3_strm1_data_mask   ;
  input                                           std__pe52__lane3_strm1_data_valid  ;

  output                                          pe52__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane4_strm0_data_mask   ;
  input                                           std__pe52__lane4_strm0_data_valid  ;

  output                                          pe52__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane4_strm1_data_mask   ;
  input                                           std__pe52__lane4_strm1_data_valid  ;

  output                                          pe52__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane5_strm0_data_mask   ;
  input                                           std__pe52__lane5_strm0_data_valid  ;

  output                                          pe52__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane5_strm1_data_mask   ;
  input                                           std__pe52__lane5_strm1_data_valid  ;

  output                                          pe52__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane6_strm0_data_mask   ;
  input                                           std__pe52__lane6_strm0_data_valid  ;

  output                                          pe52__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane6_strm1_data_mask   ;
  input                                           std__pe52__lane6_strm1_data_valid  ;

  output                                          pe52__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane7_strm0_data_mask   ;
  input                                           std__pe52__lane7_strm0_data_valid  ;

  output                                          pe52__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane7_strm1_data_mask   ;
  input                                           std__pe52__lane7_strm1_data_valid  ;

  output                                          pe52__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane8_strm0_data_mask   ;
  input                                           std__pe52__lane8_strm0_data_valid  ;

  output                                          pe52__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane8_strm1_data_mask   ;
  input                                           std__pe52__lane8_strm1_data_valid  ;

  output                                          pe52__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane9_strm0_data_mask   ;
  input                                           std__pe52__lane9_strm0_data_valid  ;

  output                                          pe52__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane9_strm1_data_mask   ;
  input                                           std__pe52__lane9_strm1_data_valid  ;

  output                                          pe52__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane10_strm0_data_mask   ;
  input                                           std__pe52__lane10_strm0_data_valid  ;

  output                                          pe52__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane10_strm1_data_mask   ;
  input                                           std__pe52__lane10_strm1_data_valid  ;

  output                                          pe52__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane11_strm0_data_mask   ;
  input                                           std__pe52__lane11_strm0_data_valid  ;

  output                                          pe52__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane11_strm1_data_mask   ;
  input                                           std__pe52__lane11_strm1_data_valid  ;

  output                                          pe52__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane12_strm0_data_mask   ;
  input                                           std__pe52__lane12_strm0_data_valid  ;

  output                                          pe52__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane12_strm1_data_mask   ;
  input                                           std__pe52__lane12_strm1_data_valid  ;

  output                                          pe52__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane13_strm0_data_mask   ;
  input                                           std__pe52__lane13_strm0_data_valid  ;

  output                                          pe52__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane13_strm1_data_mask   ;
  input                                           std__pe52__lane13_strm1_data_valid  ;

  output                                          pe52__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane14_strm0_data_mask   ;
  input                                           std__pe52__lane14_strm0_data_valid  ;

  output                                          pe52__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane14_strm1_data_mask   ;
  input                                           std__pe52__lane14_strm1_data_valid  ;

  output                                          pe52__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane15_strm0_data_mask   ;
  input                                           std__pe52__lane15_strm0_data_valid  ;

  output                                          pe52__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane15_strm1_data_mask   ;
  input                                           std__pe52__lane15_strm1_data_valid  ;

  output                                          pe52__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane16_strm0_data_mask   ;
  input                                           std__pe52__lane16_strm0_data_valid  ;

  output                                          pe52__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane16_strm1_data_mask   ;
  input                                           std__pe52__lane16_strm1_data_valid  ;

  output                                          pe52__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane17_strm0_data_mask   ;
  input                                           std__pe52__lane17_strm0_data_valid  ;

  output                                          pe52__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane17_strm1_data_mask   ;
  input                                           std__pe52__lane17_strm1_data_valid  ;

  output                                          pe52__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane18_strm0_data_mask   ;
  input                                           std__pe52__lane18_strm0_data_valid  ;

  output                                          pe52__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane18_strm1_data_mask   ;
  input                                           std__pe52__lane18_strm1_data_valid  ;

  output                                          pe52__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane19_strm0_data_mask   ;
  input                                           std__pe52__lane19_strm0_data_valid  ;

  output                                          pe52__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane19_strm1_data_mask   ;
  input                                           std__pe52__lane19_strm1_data_valid  ;

  output                                          pe52__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane20_strm0_data_mask   ;
  input                                           std__pe52__lane20_strm0_data_valid  ;

  output                                          pe52__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane20_strm1_data_mask   ;
  input                                           std__pe52__lane20_strm1_data_valid  ;

  output                                          pe52__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane21_strm0_data_mask   ;
  input                                           std__pe52__lane21_strm0_data_valid  ;

  output                                          pe52__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane21_strm1_data_mask   ;
  input                                           std__pe52__lane21_strm1_data_valid  ;

  output                                          pe52__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane22_strm0_data_mask   ;
  input                                           std__pe52__lane22_strm0_data_valid  ;

  output                                          pe52__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane22_strm1_data_mask   ;
  input                                           std__pe52__lane22_strm1_data_valid  ;

  output                                          pe52__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane23_strm0_data_mask   ;
  input                                           std__pe52__lane23_strm0_data_valid  ;

  output                                          pe52__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane23_strm1_data_mask   ;
  input                                           std__pe52__lane23_strm1_data_valid  ;

  output                                          pe52__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane24_strm0_data_mask   ;
  input                                           std__pe52__lane24_strm0_data_valid  ;

  output                                          pe52__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane24_strm1_data_mask   ;
  input                                           std__pe52__lane24_strm1_data_valid  ;

  output                                          pe52__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane25_strm0_data_mask   ;
  input                                           std__pe52__lane25_strm0_data_valid  ;

  output                                          pe52__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane25_strm1_data_mask   ;
  input                                           std__pe52__lane25_strm1_data_valid  ;

  output                                          pe52__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane26_strm0_data_mask   ;
  input                                           std__pe52__lane26_strm0_data_valid  ;

  output                                          pe52__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane26_strm1_data_mask   ;
  input                                           std__pe52__lane26_strm1_data_valid  ;

  output                                          pe52__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane27_strm0_data_mask   ;
  input                                           std__pe52__lane27_strm0_data_valid  ;

  output                                          pe52__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane27_strm1_data_mask   ;
  input                                           std__pe52__lane27_strm1_data_valid  ;

  output                                          pe52__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane28_strm0_data_mask   ;
  input                                           std__pe52__lane28_strm0_data_valid  ;

  output                                          pe52__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane28_strm1_data_mask   ;
  input                                           std__pe52__lane28_strm1_data_valid  ;

  output                                          pe52__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane29_strm0_data_mask   ;
  input                                           std__pe52__lane29_strm0_data_valid  ;

  output                                          pe52__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane29_strm1_data_mask   ;
  input                                           std__pe52__lane29_strm1_data_valid  ;

  output                                          pe52__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane30_strm0_data_mask   ;
  input                                           std__pe52__lane30_strm0_data_valid  ;

  output                                          pe52__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane30_strm1_data_mask   ;
  input                                           std__pe52__lane30_strm1_data_valid  ;

  output                                          pe52__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane31_strm0_data_mask   ;
  input                                           std__pe52__lane31_strm0_data_valid  ;

  output                                          pe52__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe52__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe52__lane31_strm1_data_mask   ;
  input                                           std__pe52__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe53__peId                ;
  input                                         sys__pe53__allSynchronized     ;
  output                                        pe53__sys__thisSynchronized    ;
  output                                        pe53__sys__ready               ;
  output                                        pe53__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe53__oob_cntl            ;
  input                                         std__pe53__oob_valid           ;
  output                                        pe53__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe53__oob_type            ;
  output                                          pe53__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane0_strm0_data_mask   ;
  input                                           std__pe53__lane0_strm0_data_valid  ;

  output                                          pe53__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane0_strm1_data_mask   ;
  input                                           std__pe53__lane0_strm1_data_valid  ;

  output                                          pe53__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane1_strm0_data_mask   ;
  input                                           std__pe53__lane1_strm0_data_valid  ;

  output                                          pe53__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane1_strm1_data_mask   ;
  input                                           std__pe53__lane1_strm1_data_valid  ;

  output                                          pe53__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane2_strm0_data_mask   ;
  input                                           std__pe53__lane2_strm0_data_valid  ;

  output                                          pe53__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane2_strm1_data_mask   ;
  input                                           std__pe53__lane2_strm1_data_valid  ;

  output                                          pe53__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane3_strm0_data_mask   ;
  input                                           std__pe53__lane3_strm0_data_valid  ;

  output                                          pe53__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane3_strm1_data_mask   ;
  input                                           std__pe53__lane3_strm1_data_valid  ;

  output                                          pe53__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane4_strm0_data_mask   ;
  input                                           std__pe53__lane4_strm0_data_valid  ;

  output                                          pe53__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane4_strm1_data_mask   ;
  input                                           std__pe53__lane4_strm1_data_valid  ;

  output                                          pe53__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane5_strm0_data_mask   ;
  input                                           std__pe53__lane5_strm0_data_valid  ;

  output                                          pe53__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane5_strm1_data_mask   ;
  input                                           std__pe53__lane5_strm1_data_valid  ;

  output                                          pe53__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane6_strm0_data_mask   ;
  input                                           std__pe53__lane6_strm0_data_valid  ;

  output                                          pe53__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane6_strm1_data_mask   ;
  input                                           std__pe53__lane6_strm1_data_valid  ;

  output                                          pe53__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane7_strm0_data_mask   ;
  input                                           std__pe53__lane7_strm0_data_valid  ;

  output                                          pe53__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane7_strm1_data_mask   ;
  input                                           std__pe53__lane7_strm1_data_valid  ;

  output                                          pe53__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane8_strm0_data_mask   ;
  input                                           std__pe53__lane8_strm0_data_valid  ;

  output                                          pe53__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane8_strm1_data_mask   ;
  input                                           std__pe53__lane8_strm1_data_valid  ;

  output                                          pe53__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane9_strm0_data_mask   ;
  input                                           std__pe53__lane9_strm0_data_valid  ;

  output                                          pe53__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane9_strm1_data_mask   ;
  input                                           std__pe53__lane9_strm1_data_valid  ;

  output                                          pe53__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane10_strm0_data_mask   ;
  input                                           std__pe53__lane10_strm0_data_valid  ;

  output                                          pe53__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane10_strm1_data_mask   ;
  input                                           std__pe53__lane10_strm1_data_valid  ;

  output                                          pe53__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane11_strm0_data_mask   ;
  input                                           std__pe53__lane11_strm0_data_valid  ;

  output                                          pe53__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane11_strm1_data_mask   ;
  input                                           std__pe53__lane11_strm1_data_valid  ;

  output                                          pe53__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane12_strm0_data_mask   ;
  input                                           std__pe53__lane12_strm0_data_valid  ;

  output                                          pe53__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane12_strm1_data_mask   ;
  input                                           std__pe53__lane12_strm1_data_valid  ;

  output                                          pe53__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane13_strm0_data_mask   ;
  input                                           std__pe53__lane13_strm0_data_valid  ;

  output                                          pe53__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane13_strm1_data_mask   ;
  input                                           std__pe53__lane13_strm1_data_valid  ;

  output                                          pe53__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane14_strm0_data_mask   ;
  input                                           std__pe53__lane14_strm0_data_valid  ;

  output                                          pe53__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane14_strm1_data_mask   ;
  input                                           std__pe53__lane14_strm1_data_valid  ;

  output                                          pe53__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane15_strm0_data_mask   ;
  input                                           std__pe53__lane15_strm0_data_valid  ;

  output                                          pe53__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane15_strm1_data_mask   ;
  input                                           std__pe53__lane15_strm1_data_valid  ;

  output                                          pe53__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane16_strm0_data_mask   ;
  input                                           std__pe53__lane16_strm0_data_valid  ;

  output                                          pe53__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane16_strm1_data_mask   ;
  input                                           std__pe53__lane16_strm1_data_valid  ;

  output                                          pe53__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane17_strm0_data_mask   ;
  input                                           std__pe53__lane17_strm0_data_valid  ;

  output                                          pe53__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane17_strm1_data_mask   ;
  input                                           std__pe53__lane17_strm1_data_valid  ;

  output                                          pe53__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane18_strm0_data_mask   ;
  input                                           std__pe53__lane18_strm0_data_valid  ;

  output                                          pe53__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane18_strm1_data_mask   ;
  input                                           std__pe53__lane18_strm1_data_valid  ;

  output                                          pe53__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane19_strm0_data_mask   ;
  input                                           std__pe53__lane19_strm0_data_valid  ;

  output                                          pe53__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane19_strm1_data_mask   ;
  input                                           std__pe53__lane19_strm1_data_valid  ;

  output                                          pe53__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane20_strm0_data_mask   ;
  input                                           std__pe53__lane20_strm0_data_valid  ;

  output                                          pe53__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane20_strm1_data_mask   ;
  input                                           std__pe53__lane20_strm1_data_valid  ;

  output                                          pe53__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane21_strm0_data_mask   ;
  input                                           std__pe53__lane21_strm0_data_valid  ;

  output                                          pe53__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane21_strm1_data_mask   ;
  input                                           std__pe53__lane21_strm1_data_valid  ;

  output                                          pe53__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane22_strm0_data_mask   ;
  input                                           std__pe53__lane22_strm0_data_valid  ;

  output                                          pe53__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane22_strm1_data_mask   ;
  input                                           std__pe53__lane22_strm1_data_valid  ;

  output                                          pe53__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane23_strm0_data_mask   ;
  input                                           std__pe53__lane23_strm0_data_valid  ;

  output                                          pe53__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane23_strm1_data_mask   ;
  input                                           std__pe53__lane23_strm1_data_valid  ;

  output                                          pe53__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane24_strm0_data_mask   ;
  input                                           std__pe53__lane24_strm0_data_valid  ;

  output                                          pe53__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane24_strm1_data_mask   ;
  input                                           std__pe53__lane24_strm1_data_valid  ;

  output                                          pe53__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane25_strm0_data_mask   ;
  input                                           std__pe53__lane25_strm0_data_valid  ;

  output                                          pe53__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane25_strm1_data_mask   ;
  input                                           std__pe53__lane25_strm1_data_valid  ;

  output                                          pe53__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane26_strm0_data_mask   ;
  input                                           std__pe53__lane26_strm0_data_valid  ;

  output                                          pe53__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane26_strm1_data_mask   ;
  input                                           std__pe53__lane26_strm1_data_valid  ;

  output                                          pe53__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane27_strm0_data_mask   ;
  input                                           std__pe53__lane27_strm0_data_valid  ;

  output                                          pe53__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane27_strm1_data_mask   ;
  input                                           std__pe53__lane27_strm1_data_valid  ;

  output                                          pe53__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane28_strm0_data_mask   ;
  input                                           std__pe53__lane28_strm0_data_valid  ;

  output                                          pe53__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane28_strm1_data_mask   ;
  input                                           std__pe53__lane28_strm1_data_valid  ;

  output                                          pe53__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane29_strm0_data_mask   ;
  input                                           std__pe53__lane29_strm0_data_valid  ;

  output                                          pe53__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane29_strm1_data_mask   ;
  input                                           std__pe53__lane29_strm1_data_valid  ;

  output                                          pe53__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane30_strm0_data_mask   ;
  input                                           std__pe53__lane30_strm0_data_valid  ;

  output                                          pe53__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane30_strm1_data_mask   ;
  input                                           std__pe53__lane30_strm1_data_valid  ;

  output                                          pe53__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane31_strm0_data_mask   ;
  input                                           std__pe53__lane31_strm0_data_valid  ;

  output                                          pe53__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe53__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe53__lane31_strm1_data_mask   ;
  input                                           std__pe53__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe54__peId                ;
  input                                         sys__pe54__allSynchronized     ;
  output                                        pe54__sys__thisSynchronized    ;
  output                                        pe54__sys__ready               ;
  output                                        pe54__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe54__oob_cntl            ;
  input                                         std__pe54__oob_valid           ;
  output                                        pe54__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe54__oob_type            ;
  output                                          pe54__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane0_strm0_data_mask   ;
  input                                           std__pe54__lane0_strm0_data_valid  ;

  output                                          pe54__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane0_strm1_data_mask   ;
  input                                           std__pe54__lane0_strm1_data_valid  ;

  output                                          pe54__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane1_strm0_data_mask   ;
  input                                           std__pe54__lane1_strm0_data_valid  ;

  output                                          pe54__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane1_strm1_data_mask   ;
  input                                           std__pe54__lane1_strm1_data_valid  ;

  output                                          pe54__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane2_strm0_data_mask   ;
  input                                           std__pe54__lane2_strm0_data_valid  ;

  output                                          pe54__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane2_strm1_data_mask   ;
  input                                           std__pe54__lane2_strm1_data_valid  ;

  output                                          pe54__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane3_strm0_data_mask   ;
  input                                           std__pe54__lane3_strm0_data_valid  ;

  output                                          pe54__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane3_strm1_data_mask   ;
  input                                           std__pe54__lane3_strm1_data_valid  ;

  output                                          pe54__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane4_strm0_data_mask   ;
  input                                           std__pe54__lane4_strm0_data_valid  ;

  output                                          pe54__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane4_strm1_data_mask   ;
  input                                           std__pe54__lane4_strm1_data_valid  ;

  output                                          pe54__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane5_strm0_data_mask   ;
  input                                           std__pe54__lane5_strm0_data_valid  ;

  output                                          pe54__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane5_strm1_data_mask   ;
  input                                           std__pe54__lane5_strm1_data_valid  ;

  output                                          pe54__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane6_strm0_data_mask   ;
  input                                           std__pe54__lane6_strm0_data_valid  ;

  output                                          pe54__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane6_strm1_data_mask   ;
  input                                           std__pe54__lane6_strm1_data_valid  ;

  output                                          pe54__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane7_strm0_data_mask   ;
  input                                           std__pe54__lane7_strm0_data_valid  ;

  output                                          pe54__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane7_strm1_data_mask   ;
  input                                           std__pe54__lane7_strm1_data_valid  ;

  output                                          pe54__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane8_strm0_data_mask   ;
  input                                           std__pe54__lane8_strm0_data_valid  ;

  output                                          pe54__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane8_strm1_data_mask   ;
  input                                           std__pe54__lane8_strm1_data_valid  ;

  output                                          pe54__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane9_strm0_data_mask   ;
  input                                           std__pe54__lane9_strm0_data_valid  ;

  output                                          pe54__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane9_strm1_data_mask   ;
  input                                           std__pe54__lane9_strm1_data_valid  ;

  output                                          pe54__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane10_strm0_data_mask   ;
  input                                           std__pe54__lane10_strm0_data_valid  ;

  output                                          pe54__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane10_strm1_data_mask   ;
  input                                           std__pe54__lane10_strm1_data_valid  ;

  output                                          pe54__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane11_strm0_data_mask   ;
  input                                           std__pe54__lane11_strm0_data_valid  ;

  output                                          pe54__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane11_strm1_data_mask   ;
  input                                           std__pe54__lane11_strm1_data_valid  ;

  output                                          pe54__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane12_strm0_data_mask   ;
  input                                           std__pe54__lane12_strm0_data_valid  ;

  output                                          pe54__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane12_strm1_data_mask   ;
  input                                           std__pe54__lane12_strm1_data_valid  ;

  output                                          pe54__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane13_strm0_data_mask   ;
  input                                           std__pe54__lane13_strm0_data_valid  ;

  output                                          pe54__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane13_strm1_data_mask   ;
  input                                           std__pe54__lane13_strm1_data_valid  ;

  output                                          pe54__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane14_strm0_data_mask   ;
  input                                           std__pe54__lane14_strm0_data_valid  ;

  output                                          pe54__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane14_strm1_data_mask   ;
  input                                           std__pe54__lane14_strm1_data_valid  ;

  output                                          pe54__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane15_strm0_data_mask   ;
  input                                           std__pe54__lane15_strm0_data_valid  ;

  output                                          pe54__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane15_strm1_data_mask   ;
  input                                           std__pe54__lane15_strm1_data_valid  ;

  output                                          pe54__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane16_strm0_data_mask   ;
  input                                           std__pe54__lane16_strm0_data_valid  ;

  output                                          pe54__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane16_strm1_data_mask   ;
  input                                           std__pe54__lane16_strm1_data_valid  ;

  output                                          pe54__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane17_strm0_data_mask   ;
  input                                           std__pe54__lane17_strm0_data_valid  ;

  output                                          pe54__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane17_strm1_data_mask   ;
  input                                           std__pe54__lane17_strm1_data_valid  ;

  output                                          pe54__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane18_strm0_data_mask   ;
  input                                           std__pe54__lane18_strm0_data_valid  ;

  output                                          pe54__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane18_strm1_data_mask   ;
  input                                           std__pe54__lane18_strm1_data_valid  ;

  output                                          pe54__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane19_strm0_data_mask   ;
  input                                           std__pe54__lane19_strm0_data_valid  ;

  output                                          pe54__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane19_strm1_data_mask   ;
  input                                           std__pe54__lane19_strm1_data_valid  ;

  output                                          pe54__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane20_strm0_data_mask   ;
  input                                           std__pe54__lane20_strm0_data_valid  ;

  output                                          pe54__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane20_strm1_data_mask   ;
  input                                           std__pe54__lane20_strm1_data_valid  ;

  output                                          pe54__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane21_strm0_data_mask   ;
  input                                           std__pe54__lane21_strm0_data_valid  ;

  output                                          pe54__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane21_strm1_data_mask   ;
  input                                           std__pe54__lane21_strm1_data_valid  ;

  output                                          pe54__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane22_strm0_data_mask   ;
  input                                           std__pe54__lane22_strm0_data_valid  ;

  output                                          pe54__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane22_strm1_data_mask   ;
  input                                           std__pe54__lane22_strm1_data_valid  ;

  output                                          pe54__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane23_strm0_data_mask   ;
  input                                           std__pe54__lane23_strm0_data_valid  ;

  output                                          pe54__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane23_strm1_data_mask   ;
  input                                           std__pe54__lane23_strm1_data_valid  ;

  output                                          pe54__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane24_strm0_data_mask   ;
  input                                           std__pe54__lane24_strm0_data_valid  ;

  output                                          pe54__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane24_strm1_data_mask   ;
  input                                           std__pe54__lane24_strm1_data_valid  ;

  output                                          pe54__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane25_strm0_data_mask   ;
  input                                           std__pe54__lane25_strm0_data_valid  ;

  output                                          pe54__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane25_strm1_data_mask   ;
  input                                           std__pe54__lane25_strm1_data_valid  ;

  output                                          pe54__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane26_strm0_data_mask   ;
  input                                           std__pe54__lane26_strm0_data_valid  ;

  output                                          pe54__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane26_strm1_data_mask   ;
  input                                           std__pe54__lane26_strm1_data_valid  ;

  output                                          pe54__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane27_strm0_data_mask   ;
  input                                           std__pe54__lane27_strm0_data_valid  ;

  output                                          pe54__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane27_strm1_data_mask   ;
  input                                           std__pe54__lane27_strm1_data_valid  ;

  output                                          pe54__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane28_strm0_data_mask   ;
  input                                           std__pe54__lane28_strm0_data_valid  ;

  output                                          pe54__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane28_strm1_data_mask   ;
  input                                           std__pe54__lane28_strm1_data_valid  ;

  output                                          pe54__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane29_strm0_data_mask   ;
  input                                           std__pe54__lane29_strm0_data_valid  ;

  output                                          pe54__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane29_strm1_data_mask   ;
  input                                           std__pe54__lane29_strm1_data_valid  ;

  output                                          pe54__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane30_strm0_data_mask   ;
  input                                           std__pe54__lane30_strm0_data_valid  ;

  output                                          pe54__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane30_strm1_data_mask   ;
  input                                           std__pe54__lane30_strm1_data_valid  ;

  output                                          pe54__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane31_strm0_data_mask   ;
  input                                           std__pe54__lane31_strm0_data_valid  ;

  output                                          pe54__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe54__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe54__lane31_strm1_data_mask   ;
  input                                           std__pe54__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe55__peId                ;
  input                                         sys__pe55__allSynchronized     ;
  output                                        pe55__sys__thisSynchronized    ;
  output                                        pe55__sys__ready               ;
  output                                        pe55__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe55__oob_cntl            ;
  input                                         std__pe55__oob_valid           ;
  output                                        pe55__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe55__oob_type            ;
  output                                          pe55__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane0_strm0_data_mask   ;
  input                                           std__pe55__lane0_strm0_data_valid  ;

  output                                          pe55__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane0_strm1_data_mask   ;
  input                                           std__pe55__lane0_strm1_data_valid  ;

  output                                          pe55__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane1_strm0_data_mask   ;
  input                                           std__pe55__lane1_strm0_data_valid  ;

  output                                          pe55__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane1_strm1_data_mask   ;
  input                                           std__pe55__lane1_strm1_data_valid  ;

  output                                          pe55__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane2_strm0_data_mask   ;
  input                                           std__pe55__lane2_strm0_data_valid  ;

  output                                          pe55__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane2_strm1_data_mask   ;
  input                                           std__pe55__lane2_strm1_data_valid  ;

  output                                          pe55__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane3_strm0_data_mask   ;
  input                                           std__pe55__lane3_strm0_data_valid  ;

  output                                          pe55__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane3_strm1_data_mask   ;
  input                                           std__pe55__lane3_strm1_data_valid  ;

  output                                          pe55__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane4_strm0_data_mask   ;
  input                                           std__pe55__lane4_strm0_data_valid  ;

  output                                          pe55__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane4_strm1_data_mask   ;
  input                                           std__pe55__lane4_strm1_data_valid  ;

  output                                          pe55__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane5_strm0_data_mask   ;
  input                                           std__pe55__lane5_strm0_data_valid  ;

  output                                          pe55__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane5_strm1_data_mask   ;
  input                                           std__pe55__lane5_strm1_data_valid  ;

  output                                          pe55__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane6_strm0_data_mask   ;
  input                                           std__pe55__lane6_strm0_data_valid  ;

  output                                          pe55__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane6_strm1_data_mask   ;
  input                                           std__pe55__lane6_strm1_data_valid  ;

  output                                          pe55__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane7_strm0_data_mask   ;
  input                                           std__pe55__lane7_strm0_data_valid  ;

  output                                          pe55__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane7_strm1_data_mask   ;
  input                                           std__pe55__lane7_strm1_data_valid  ;

  output                                          pe55__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane8_strm0_data_mask   ;
  input                                           std__pe55__lane8_strm0_data_valid  ;

  output                                          pe55__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane8_strm1_data_mask   ;
  input                                           std__pe55__lane8_strm1_data_valid  ;

  output                                          pe55__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane9_strm0_data_mask   ;
  input                                           std__pe55__lane9_strm0_data_valid  ;

  output                                          pe55__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane9_strm1_data_mask   ;
  input                                           std__pe55__lane9_strm1_data_valid  ;

  output                                          pe55__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane10_strm0_data_mask   ;
  input                                           std__pe55__lane10_strm0_data_valid  ;

  output                                          pe55__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane10_strm1_data_mask   ;
  input                                           std__pe55__lane10_strm1_data_valid  ;

  output                                          pe55__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane11_strm0_data_mask   ;
  input                                           std__pe55__lane11_strm0_data_valid  ;

  output                                          pe55__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane11_strm1_data_mask   ;
  input                                           std__pe55__lane11_strm1_data_valid  ;

  output                                          pe55__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane12_strm0_data_mask   ;
  input                                           std__pe55__lane12_strm0_data_valid  ;

  output                                          pe55__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane12_strm1_data_mask   ;
  input                                           std__pe55__lane12_strm1_data_valid  ;

  output                                          pe55__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane13_strm0_data_mask   ;
  input                                           std__pe55__lane13_strm0_data_valid  ;

  output                                          pe55__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane13_strm1_data_mask   ;
  input                                           std__pe55__lane13_strm1_data_valid  ;

  output                                          pe55__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane14_strm0_data_mask   ;
  input                                           std__pe55__lane14_strm0_data_valid  ;

  output                                          pe55__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane14_strm1_data_mask   ;
  input                                           std__pe55__lane14_strm1_data_valid  ;

  output                                          pe55__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane15_strm0_data_mask   ;
  input                                           std__pe55__lane15_strm0_data_valid  ;

  output                                          pe55__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane15_strm1_data_mask   ;
  input                                           std__pe55__lane15_strm1_data_valid  ;

  output                                          pe55__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane16_strm0_data_mask   ;
  input                                           std__pe55__lane16_strm0_data_valid  ;

  output                                          pe55__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane16_strm1_data_mask   ;
  input                                           std__pe55__lane16_strm1_data_valid  ;

  output                                          pe55__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane17_strm0_data_mask   ;
  input                                           std__pe55__lane17_strm0_data_valid  ;

  output                                          pe55__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane17_strm1_data_mask   ;
  input                                           std__pe55__lane17_strm1_data_valid  ;

  output                                          pe55__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane18_strm0_data_mask   ;
  input                                           std__pe55__lane18_strm0_data_valid  ;

  output                                          pe55__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane18_strm1_data_mask   ;
  input                                           std__pe55__lane18_strm1_data_valid  ;

  output                                          pe55__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane19_strm0_data_mask   ;
  input                                           std__pe55__lane19_strm0_data_valid  ;

  output                                          pe55__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane19_strm1_data_mask   ;
  input                                           std__pe55__lane19_strm1_data_valid  ;

  output                                          pe55__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane20_strm0_data_mask   ;
  input                                           std__pe55__lane20_strm0_data_valid  ;

  output                                          pe55__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane20_strm1_data_mask   ;
  input                                           std__pe55__lane20_strm1_data_valid  ;

  output                                          pe55__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane21_strm0_data_mask   ;
  input                                           std__pe55__lane21_strm0_data_valid  ;

  output                                          pe55__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane21_strm1_data_mask   ;
  input                                           std__pe55__lane21_strm1_data_valid  ;

  output                                          pe55__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane22_strm0_data_mask   ;
  input                                           std__pe55__lane22_strm0_data_valid  ;

  output                                          pe55__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane22_strm1_data_mask   ;
  input                                           std__pe55__lane22_strm1_data_valid  ;

  output                                          pe55__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane23_strm0_data_mask   ;
  input                                           std__pe55__lane23_strm0_data_valid  ;

  output                                          pe55__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane23_strm1_data_mask   ;
  input                                           std__pe55__lane23_strm1_data_valid  ;

  output                                          pe55__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane24_strm0_data_mask   ;
  input                                           std__pe55__lane24_strm0_data_valid  ;

  output                                          pe55__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane24_strm1_data_mask   ;
  input                                           std__pe55__lane24_strm1_data_valid  ;

  output                                          pe55__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane25_strm0_data_mask   ;
  input                                           std__pe55__lane25_strm0_data_valid  ;

  output                                          pe55__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane25_strm1_data_mask   ;
  input                                           std__pe55__lane25_strm1_data_valid  ;

  output                                          pe55__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane26_strm0_data_mask   ;
  input                                           std__pe55__lane26_strm0_data_valid  ;

  output                                          pe55__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane26_strm1_data_mask   ;
  input                                           std__pe55__lane26_strm1_data_valid  ;

  output                                          pe55__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane27_strm0_data_mask   ;
  input                                           std__pe55__lane27_strm0_data_valid  ;

  output                                          pe55__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane27_strm1_data_mask   ;
  input                                           std__pe55__lane27_strm1_data_valid  ;

  output                                          pe55__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane28_strm0_data_mask   ;
  input                                           std__pe55__lane28_strm0_data_valid  ;

  output                                          pe55__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane28_strm1_data_mask   ;
  input                                           std__pe55__lane28_strm1_data_valid  ;

  output                                          pe55__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane29_strm0_data_mask   ;
  input                                           std__pe55__lane29_strm0_data_valid  ;

  output                                          pe55__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane29_strm1_data_mask   ;
  input                                           std__pe55__lane29_strm1_data_valid  ;

  output                                          pe55__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane30_strm0_data_mask   ;
  input                                           std__pe55__lane30_strm0_data_valid  ;

  output                                          pe55__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane30_strm1_data_mask   ;
  input                                           std__pe55__lane30_strm1_data_valid  ;

  output                                          pe55__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane31_strm0_data_mask   ;
  input                                           std__pe55__lane31_strm0_data_valid  ;

  output                                          pe55__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe55__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe55__lane31_strm1_data_mask   ;
  input                                           std__pe55__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe56__peId                ;
  input                                         sys__pe56__allSynchronized     ;
  output                                        pe56__sys__thisSynchronized    ;
  output                                        pe56__sys__ready               ;
  output                                        pe56__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe56__oob_cntl            ;
  input                                         std__pe56__oob_valid           ;
  output                                        pe56__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe56__oob_type            ;
  output                                          pe56__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane0_strm0_data_mask   ;
  input                                           std__pe56__lane0_strm0_data_valid  ;

  output                                          pe56__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane0_strm1_data_mask   ;
  input                                           std__pe56__lane0_strm1_data_valid  ;

  output                                          pe56__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane1_strm0_data_mask   ;
  input                                           std__pe56__lane1_strm0_data_valid  ;

  output                                          pe56__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane1_strm1_data_mask   ;
  input                                           std__pe56__lane1_strm1_data_valid  ;

  output                                          pe56__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane2_strm0_data_mask   ;
  input                                           std__pe56__lane2_strm0_data_valid  ;

  output                                          pe56__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane2_strm1_data_mask   ;
  input                                           std__pe56__lane2_strm1_data_valid  ;

  output                                          pe56__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane3_strm0_data_mask   ;
  input                                           std__pe56__lane3_strm0_data_valid  ;

  output                                          pe56__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane3_strm1_data_mask   ;
  input                                           std__pe56__lane3_strm1_data_valid  ;

  output                                          pe56__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane4_strm0_data_mask   ;
  input                                           std__pe56__lane4_strm0_data_valid  ;

  output                                          pe56__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane4_strm1_data_mask   ;
  input                                           std__pe56__lane4_strm1_data_valid  ;

  output                                          pe56__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane5_strm0_data_mask   ;
  input                                           std__pe56__lane5_strm0_data_valid  ;

  output                                          pe56__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane5_strm1_data_mask   ;
  input                                           std__pe56__lane5_strm1_data_valid  ;

  output                                          pe56__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane6_strm0_data_mask   ;
  input                                           std__pe56__lane6_strm0_data_valid  ;

  output                                          pe56__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane6_strm1_data_mask   ;
  input                                           std__pe56__lane6_strm1_data_valid  ;

  output                                          pe56__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane7_strm0_data_mask   ;
  input                                           std__pe56__lane7_strm0_data_valid  ;

  output                                          pe56__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane7_strm1_data_mask   ;
  input                                           std__pe56__lane7_strm1_data_valid  ;

  output                                          pe56__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane8_strm0_data_mask   ;
  input                                           std__pe56__lane8_strm0_data_valid  ;

  output                                          pe56__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane8_strm1_data_mask   ;
  input                                           std__pe56__lane8_strm1_data_valid  ;

  output                                          pe56__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane9_strm0_data_mask   ;
  input                                           std__pe56__lane9_strm0_data_valid  ;

  output                                          pe56__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane9_strm1_data_mask   ;
  input                                           std__pe56__lane9_strm1_data_valid  ;

  output                                          pe56__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane10_strm0_data_mask   ;
  input                                           std__pe56__lane10_strm0_data_valid  ;

  output                                          pe56__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane10_strm1_data_mask   ;
  input                                           std__pe56__lane10_strm1_data_valid  ;

  output                                          pe56__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane11_strm0_data_mask   ;
  input                                           std__pe56__lane11_strm0_data_valid  ;

  output                                          pe56__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane11_strm1_data_mask   ;
  input                                           std__pe56__lane11_strm1_data_valid  ;

  output                                          pe56__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane12_strm0_data_mask   ;
  input                                           std__pe56__lane12_strm0_data_valid  ;

  output                                          pe56__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane12_strm1_data_mask   ;
  input                                           std__pe56__lane12_strm1_data_valid  ;

  output                                          pe56__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane13_strm0_data_mask   ;
  input                                           std__pe56__lane13_strm0_data_valid  ;

  output                                          pe56__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane13_strm1_data_mask   ;
  input                                           std__pe56__lane13_strm1_data_valid  ;

  output                                          pe56__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane14_strm0_data_mask   ;
  input                                           std__pe56__lane14_strm0_data_valid  ;

  output                                          pe56__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane14_strm1_data_mask   ;
  input                                           std__pe56__lane14_strm1_data_valid  ;

  output                                          pe56__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane15_strm0_data_mask   ;
  input                                           std__pe56__lane15_strm0_data_valid  ;

  output                                          pe56__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane15_strm1_data_mask   ;
  input                                           std__pe56__lane15_strm1_data_valid  ;

  output                                          pe56__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane16_strm0_data_mask   ;
  input                                           std__pe56__lane16_strm0_data_valid  ;

  output                                          pe56__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane16_strm1_data_mask   ;
  input                                           std__pe56__lane16_strm1_data_valid  ;

  output                                          pe56__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane17_strm0_data_mask   ;
  input                                           std__pe56__lane17_strm0_data_valid  ;

  output                                          pe56__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane17_strm1_data_mask   ;
  input                                           std__pe56__lane17_strm1_data_valid  ;

  output                                          pe56__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane18_strm0_data_mask   ;
  input                                           std__pe56__lane18_strm0_data_valid  ;

  output                                          pe56__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane18_strm1_data_mask   ;
  input                                           std__pe56__lane18_strm1_data_valid  ;

  output                                          pe56__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane19_strm0_data_mask   ;
  input                                           std__pe56__lane19_strm0_data_valid  ;

  output                                          pe56__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane19_strm1_data_mask   ;
  input                                           std__pe56__lane19_strm1_data_valid  ;

  output                                          pe56__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane20_strm0_data_mask   ;
  input                                           std__pe56__lane20_strm0_data_valid  ;

  output                                          pe56__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane20_strm1_data_mask   ;
  input                                           std__pe56__lane20_strm1_data_valid  ;

  output                                          pe56__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane21_strm0_data_mask   ;
  input                                           std__pe56__lane21_strm0_data_valid  ;

  output                                          pe56__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane21_strm1_data_mask   ;
  input                                           std__pe56__lane21_strm1_data_valid  ;

  output                                          pe56__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane22_strm0_data_mask   ;
  input                                           std__pe56__lane22_strm0_data_valid  ;

  output                                          pe56__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane22_strm1_data_mask   ;
  input                                           std__pe56__lane22_strm1_data_valid  ;

  output                                          pe56__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane23_strm0_data_mask   ;
  input                                           std__pe56__lane23_strm0_data_valid  ;

  output                                          pe56__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane23_strm1_data_mask   ;
  input                                           std__pe56__lane23_strm1_data_valid  ;

  output                                          pe56__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane24_strm0_data_mask   ;
  input                                           std__pe56__lane24_strm0_data_valid  ;

  output                                          pe56__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane24_strm1_data_mask   ;
  input                                           std__pe56__lane24_strm1_data_valid  ;

  output                                          pe56__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane25_strm0_data_mask   ;
  input                                           std__pe56__lane25_strm0_data_valid  ;

  output                                          pe56__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane25_strm1_data_mask   ;
  input                                           std__pe56__lane25_strm1_data_valid  ;

  output                                          pe56__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane26_strm0_data_mask   ;
  input                                           std__pe56__lane26_strm0_data_valid  ;

  output                                          pe56__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane26_strm1_data_mask   ;
  input                                           std__pe56__lane26_strm1_data_valid  ;

  output                                          pe56__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane27_strm0_data_mask   ;
  input                                           std__pe56__lane27_strm0_data_valid  ;

  output                                          pe56__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane27_strm1_data_mask   ;
  input                                           std__pe56__lane27_strm1_data_valid  ;

  output                                          pe56__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane28_strm0_data_mask   ;
  input                                           std__pe56__lane28_strm0_data_valid  ;

  output                                          pe56__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane28_strm1_data_mask   ;
  input                                           std__pe56__lane28_strm1_data_valid  ;

  output                                          pe56__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane29_strm0_data_mask   ;
  input                                           std__pe56__lane29_strm0_data_valid  ;

  output                                          pe56__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane29_strm1_data_mask   ;
  input                                           std__pe56__lane29_strm1_data_valid  ;

  output                                          pe56__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane30_strm0_data_mask   ;
  input                                           std__pe56__lane30_strm0_data_valid  ;

  output                                          pe56__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane30_strm1_data_mask   ;
  input                                           std__pe56__lane30_strm1_data_valid  ;

  output                                          pe56__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane31_strm0_data_mask   ;
  input                                           std__pe56__lane31_strm0_data_valid  ;

  output                                          pe56__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe56__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe56__lane31_strm1_data_mask   ;
  input                                           std__pe56__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe57__peId                ;
  input                                         sys__pe57__allSynchronized     ;
  output                                        pe57__sys__thisSynchronized    ;
  output                                        pe57__sys__ready               ;
  output                                        pe57__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe57__oob_cntl            ;
  input                                         std__pe57__oob_valid           ;
  output                                        pe57__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe57__oob_type            ;
  output                                          pe57__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane0_strm0_data_mask   ;
  input                                           std__pe57__lane0_strm0_data_valid  ;

  output                                          pe57__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane0_strm1_data_mask   ;
  input                                           std__pe57__lane0_strm1_data_valid  ;

  output                                          pe57__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane1_strm0_data_mask   ;
  input                                           std__pe57__lane1_strm0_data_valid  ;

  output                                          pe57__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane1_strm1_data_mask   ;
  input                                           std__pe57__lane1_strm1_data_valid  ;

  output                                          pe57__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane2_strm0_data_mask   ;
  input                                           std__pe57__lane2_strm0_data_valid  ;

  output                                          pe57__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane2_strm1_data_mask   ;
  input                                           std__pe57__lane2_strm1_data_valid  ;

  output                                          pe57__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane3_strm0_data_mask   ;
  input                                           std__pe57__lane3_strm0_data_valid  ;

  output                                          pe57__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane3_strm1_data_mask   ;
  input                                           std__pe57__lane3_strm1_data_valid  ;

  output                                          pe57__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane4_strm0_data_mask   ;
  input                                           std__pe57__lane4_strm0_data_valid  ;

  output                                          pe57__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane4_strm1_data_mask   ;
  input                                           std__pe57__lane4_strm1_data_valid  ;

  output                                          pe57__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane5_strm0_data_mask   ;
  input                                           std__pe57__lane5_strm0_data_valid  ;

  output                                          pe57__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane5_strm1_data_mask   ;
  input                                           std__pe57__lane5_strm1_data_valid  ;

  output                                          pe57__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane6_strm0_data_mask   ;
  input                                           std__pe57__lane6_strm0_data_valid  ;

  output                                          pe57__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane6_strm1_data_mask   ;
  input                                           std__pe57__lane6_strm1_data_valid  ;

  output                                          pe57__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane7_strm0_data_mask   ;
  input                                           std__pe57__lane7_strm0_data_valid  ;

  output                                          pe57__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane7_strm1_data_mask   ;
  input                                           std__pe57__lane7_strm1_data_valid  ;

  output                                          pe57__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane8_strm0_data_mask   ;
  input                                           std__pe57__lane8_strm0_data_valid  ;

  output                                          pe57__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane8_strm1_data_mask   ;
  input                                           std__pe57__lane8_strm1_data_valid  ;

  output                                          pe57__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane9_strm0_data_mask   ;
  input                                           std__pe57__lane9_strm0_data_valid  ;

  output                                          pe57__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane9_strm1_data_mask   ;
  input                                           std__pe57__lane9_strm1_data_valid  ;

  output                                          pe57__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane10_strm0_data_mask   ;
  input                                           std__pe57__lane10_strm0_data_valid  ;

  output                                          pe57__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane10_strm1_data_mask   ;
  input                                           std__pe57__lane10_strm1_data_valid  ;

  output                                          pe57__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane11_strm0_data_mask   ;
  input                                           std__pe57__lane11_strm0_data_valid  ;

  output                                          pe57__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane11_strm1_data_mask   ;
  input                                           std__pe57__lane11_strm1_data_valid  ;

  output                                          pe57__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane12_strm0_data_mask   ;
  input                                           std__pe57__lane12_strm0_data_valid  ;

  output                                          pe57__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane12_strm1_data_mask   ;
  input                                           std__pe57__lane12_strm1_data_valid  ;

  output                                          pe57__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane13_strm0_data_mask   ;
  input                                           std__pe57__lane13_strm0_data_valid  ;

  output                                          pe57__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane13_strm1_data_mask   ;
  input                                           std__pe57__lane13_strm1_data_valid  ;

  output                                          pe57__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane14_strm0_data_mask   ;
  input                                           std__pe57__lane14_strm0_data_valid  ;

  output                                          pe57__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane14_strm1_data_mask   ;
  input                                           std__pe57__lane14_strm1_data_valid  ;

  output                                          pe57__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane15_strm0_data_mask   ;
  input                                           std__pe57__lane15_strm0_data_valid  ;

  output                                          pe57__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane15_strm1_data_mask   ;
  input                                           std__pe57__lane15_strm1_data_valid  ;

  output                                          pe57__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane16_strm0_data_mask   ;
  input                                           std__pe57__lane16_strm0_data_valid  ;

  output                                          pe57__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane16_strm1_data_mask   ;
  input                                           std__pe57__lane16_strm1_data_valid  ;

  output                                          pe57__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane17_strm0_data_mask   ;
  input                                           std__pe57__lane17_strm0_data_valid  ;

  output                                          pe57__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane17_strm1_data_mask   ;
  input                                           std__pe57__lane17_strm1_data_valid  ;

  output                                          pe57__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane18_strm0_data_mask   ;
  input                                           std__pe57__lane18_strm0_data_valid  ;

  output                                          pe57__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane18_strm1_data_mask   ;
  input                                           std__pe57__lane18_strm1_data_valid  ;

  output                                          pe57__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane19_strm0_data_mask   ;
  input                                           std__pe57__lane19_strm0_data_valid  ;

  output                                          pe57__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane19_strm1_data_mask   ;
  input                                           std__pe57__lane19_strm1_data_valid  ;

  output                                          pe57__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane20_strm0_data_mask   ;
  input                                           std__pe57__lane20_strm0_data_valid  ;

  output                                          pe57__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane20_strm1_data_mask   ;
  input                                           std__pe57__lane20_strm1_data_valid  ;

  output                                          pe57__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane21_strm0_data_mask   ;
  input                                           std__pe57__lane21_strm0_data_valid  ;

  output                                          pe57__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane21_strm1_data_mask   ;
  input                                           std__pe57__lane21_strm1_data_valid  ;

  output                                          pe57__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane22_strm0_data_mask   ;
  input                                           std__pe57__lane22_strm0_data_valid  ;

  output                                          pe57__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane22_strm1_data_mask   ;
  input                                           std__pe57__lane22_strm1_data_valid  ;

  output                                          pe57__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane23_strm0_data_mask   ;
  input                                           std__pe57__lane23_strm0_data_valid  ;

  output                                          pe57__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane23_strm1_data_mask   ;
  input                                           std__pe57__lane23_strm1_data_valid  ;

  output                                          pe57__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane24_strm0_data_mask   ;
  input                                           std__pe57__lane24_strm0_data_valid  ;

  output                                          pe57__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane24_strm1_data_mask   ;
  input                                           std__pe57__lane24_strm1_data_valid  ;

  output                                          pe57__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane25_strm0_data_mask   ;
  input                                           std__pe57__lane25_strm0_data_valid  ;

  output                                          pe57__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane25_strm1_data_mask   ;
  input                                           std__pe57__lane25_strm1_data_valid  ;

  output                                          pe57__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane26_strm0_data_mask   ;
  input                                           std__pe57__lane26_strm0_data_valid  ;

  output                                          pe57__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane26_strm1_data_mask   ;
  input                                           std__pe57__lane26_strm1_data_valid  ;

  output                                          pe57__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane27_strm0_data_mask   ;
  input                                           std__pe57__lane27_strm0_data_valid  ;

  output                                          pe57__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane27_strm1_data_mask   ;
  input                                           std__pe57__lane27_strm1_data_valid  ;

  output                                          pe57__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane28_strm0_data_mask   ;
  input                                           std__pe57__lane28_strm0_data_valid  ;

  output                                          pe57__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane28_strm1_data_mask   ;
  input                                           std__pe57__lane28_strm1_data_valid  ;

  output                                          pe57__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane29_strm0_data_mask   ;
  input                                           std__pe57__lane29_strm0_data_valid  ;

  output                                          pe57__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane29_strm1_data_mask   ;
  input                                           std__pe57__lane29_strm1_data_valid  ;

  output                                          pe57__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane30_strm0_data_mask   ;
  input                                           std__pe57__lane30_strm0_data_valid  ;

  output                                          pe57__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane30_strm1_data_mask   ;
  input                                           std__pe57__lane30_strm1_data_valid  ;

  output                                          pe57__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane31_strm0_data_mask   ;
  input                                           std__pe57__lane31_strm0_data_valid  ;

  output                                          pe57__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe57__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe57__lane31_strm1_data_mask   ;
  input                                           std__pe57__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe58__peId                ;
  input                                         sys__pe58__allSynchronized     ;
  output                                        pe58__sys__thisSynchronized    ;
  output                                        pe58__sys__ready               ;
  output                                        pe58__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe58__oob_cntl            ;
  input                                         std__pe58__oob_valid           ;
  output                                        pe58__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe58__oob_type            ;
  output                                          pe58__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane0_strm0_data_mask   ;
  input                                           std__pe58__lane0_strm0_data_valid  ;

  output                                          pe58__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane0_strm1_data_mask   ;
  input                                           std__pe58__lane0_strm1_data_valid  ;

  output                                          pe58__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane1_strm0_data_mask   ;
  input                                           std__pe58__lane1_strm0_data_valid  ;

  output                                          pe58__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane1_strm1_data_mask   ;
  input                                           std__pe58__lane1_strm1_data_valid  ;

  output                                          pe58__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane2_strm0_data_mask   ;
  input                                           std__pe58__lane2_strm0_data_valid  ;

  output                                          pe58__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane2_strm1_data_mask   ;
  input                                           std__pe58__lane2_strm1_data_valid  ;

  output                                          pe58__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane3_strm0_data_mask   ;
  input                                           std__pe58__lane3_strm0_data_valid  ;

  output                                          pe58__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane3_strm1_data_mask   ;
  input                                           std__pe58__lane3_strm1_data_valid  ;

  output                                          pe58__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane4_strm0_data_mask   ;
  input                                           std__pe58__lane4_strm0_data_valid  ;

  output                                          pe58__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane4_strm1_data_mask   ;
  input                                           std__pe58__lane4_strm1_data_valid  ;

  output                                          pe58__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane5_strm0_data_mask   ;
  input                                           std__pe58__lane5_strm0_data_valid  ;

  output                                          pe58__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane5_strm1_data_mask   ;
  input                                           std__pe58__lane5_strm1_data_valid  ;

  output                                          pe58__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane6_strm0_data_mask   ;
  input                                           std__pe58__lane6_strm0_data_valid  ;

  output                                          pe58__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane6_strm1_data_mask   ;
  input                                           std__pe58__lane6_strm1_data_valid  ;

  output                                          pe58__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane7_strm0_data_mask   ;
  input                                           std__pe58__lane7_strm0_data_valid  ;

  output                                          pe58__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane7_strm1_data_mask   ;
  input                                           std__pe58__lane7_strm1_data_valid  ;

  output                                          pe58__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane8_strm0_data_mask   ;
  input                                           std__pe58__lane8_strm0_data_valid  ;

  output                                          pe58__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane8_strm1_data_mask   ;
  input                                           std__pe58__lane8_strm1_data_valid  ;

  output                                          pe58__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane9_strm0_data_mask   ;
  input                                           std__pe58__lane9_strm0_data_valid  ;

  output                                          pe58__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane9_strm1_data_mask   ;
  input                                           std__pe58__lane9_strm1_data_valid  ;

  output                                          pe58__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane10_strm0_data_mask   ;
  input                                           std__pe58__lane10_strm0_data_valid  ;

  output                                          pe58__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane10_strm1_data_mask   ;
  input                                           std__pe58__lane10_strm1_data_valid  ;

  output                                          pe58__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane11_strm0_data_mask   ;
  input                                           std__pe58__lane11_strm0_data_valid  ;

  output                                          pe58__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane11_strm1_data_mask   ;
  input                                           std__pe58__lane11_strm1_data_valid  ;

  output                                          pe58__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane12_strm0_data_mask   ;
  input                                           std__pe58__lane12_strm0_data_valid  ;

  output                                          pe58__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane12_strm1_data_mask   ;
  input                                           std__pe58__lane12_strm1_data_valid  ;

  output                                          pe58__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane13_strm0_data_mask   ;
  input                                           std__pe58__lane13_strm0_data_valid  ;

  output                                          pe58__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane13_strm1_data_mask   ;
  input                                           std__pe58__lane13_strm1_data_valid  ;

  output                                          pe58__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane14_strm0_data_mask   ;
  input                                           std__pe58__lane14_strm0_data_valid  ;

  output                                          pe58__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane14_strm1_data_mask   ;
  input                                           std__pe58__lane14_strm1_data_valid  ;

  output                                          pe58__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane15_strm0_data_mask   ;
  input                                           std__pe58__lane15_strm0_data_valid  ;

  output                                          pe58__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane15_strm1_data_mask   ;
  input                                           std__pe58__lane15_strm1_data_valid  ;

  output                                          pe58__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane16_strm0_data_mask   ;
  input                                           std__pe58__lane16_strm0_data_valid  ;

  output                                          pe58__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane16_strm1_data_mask   ;
  input                                           std__pe58__lane16_strm1_data_valid  ;

  output                                          pe58__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane17_strm0_data_mask   ;
  input                                           std__pe58__lane17_strm0_data_valid  ;

  output                                          pe58__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane17_strm1_data_mask   ;
  input                                           std__pe58__lane17_strm1_data_valid  ;

  output                                          pe58__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane18_strm0_data_mask   ;
  input                                           std__pe58__lane18_strm0_data_valid  ;

  output                                          pe58__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane18_strm1_data_mask   ;
  input                                           std__pe58__lane18_strm1_data_valid  ;

  output                                          pe58__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane19_strm0_data_mask   ;
  input                                           std__pe58__lane19_strm0_data_valid  ;

  output                                          pe58__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane19_strm1_data_mask   ;
  input                                           std__pe58__lane19_strm1_data_valid  ;

  output                                          pe58__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane20_strm0_data_mask   ;
  input                                           std__pe58__lane20_strm0_data_valid  ;

  output                                          pe58__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane20_strm1_data_mask   ;
  input                                           std__pe58__lane20_strm1_data_valid  ;

  output                                          pe58__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane21_strm0_data_mask   ;
  input                                           std__pe58__lane21_strm0_data_valid  ;

  output                                          pe58__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane21_strm1_data_mask   ;
  input                                           std__pe58__lane21_strm1_data_valid  ;

  output                                          pe58__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane22_strm0_data_mask   ;
  input                                           std__pe58__lane22_strm0_data_valid  ;

  output                                          pe58__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane22_strm1_data_mask   ;
  input                                           std__pe58__lane22_strm1_data_valid  ;

  output                                          pe58__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane23_strm0_data_mask   ;
  input                                           std__pe58__lane23_strm0_data_valid  ;

  output                                          pe58__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane23_strm1_data_mask   ;
  input                                           std__pe58__lane23_strm1_data_valid  ;

  output                                          pe58__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane24_strm0_data_mask   ;
  input                                           std__pe58__lane24_strm0_data_valid  ;

  output                                          pe58__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane24_strm1_data_mask   ;
  input                                           std__pe58__lane24_strm1_data_valid  ;

  output                                          pe58__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane25_strm0_data_mask   ;
  input                                           std__pe58__lane25_strm0_data_valid  ;

  output                                          pe58__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane25_strm1_data_mask   ;
  input                                           std__pe58__lane25_strm1_data_valid  ;

  output                                          pe58__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane26_strm0_data_mask   ;
  input                                           std__pe58__lane26_strm0_data_valid  ;

  output                                          pe58__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane26_strm1_data_mask   ;
  input                                           std__pe58__lane26_strm1_data_valid  ;

  output                                          pe58__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane27_strm0_data_mask   ;
  input                                           std__pe58__lane27_strm0_data_valid  ;

  output                                          pe58__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane27_strm1_data_mask   ;
  input                                           std__pe58__lane27_strm1_data_valid  ;

  output                                          pe58__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane28_strm0_data_mask   ;
  input                                           std__pe58__lane28_strm0_data_valid  ;

  output                                          pe58__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane28_strm1_data_mask   ;
  input                                           std__pe58__lane28_strm1_data_valid  ;

  output                                          pe58__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane29_strm0_data_mask   ;
  input                                           std__pe58__lane29_strm0_data_valid  ;

  output                                          pe58__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane29_strm1_data_mask   ;
  input                                           std__pe58__lane29_strm1_data_valid  ;

  output                                          pe58__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane30_strm0_data_mask   ;
  input                                           std__pe58__lane30_strm0_data_valid  ;

  output                                          pe58__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane30_strm1_data_mask   ;
  input                                           std__pe58__lane30_strm1_data_valid  ;

  output                                          pe58__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane31_strm0_data_mask   ;
  input                                           std__pe58__lane31_strm0_data_valid  ;

  output                                          pe58__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe58__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe58__lane31_strm1_data_mask   ;
  input                                           std__pe58__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe59__peId                ;
  input                                         sys__pe59__allSynchronized     ;
  output                                        pe59__sys__thisSynchronized    ;
  output                                        pe59__sys__ready               ;
  output                                        pe59__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe59__oob_cntl            ;
  input                                         std__pe59__oob_valid           ;
  output                                        pe59__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe59__oob_type            ;
  output                                          pe59__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane0_strm0_data_mask   ;
  input                                           std__pe59__lane0_strm0_data_valid  ;

  output                                          pe59__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane0_strm1_data_mask   ;
  input                                           std__pe59__lane0_strm1_data_valid  ;

  output                                          pe59__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane1_strm0_data_mask   ;
  input                                           std__pe59__lane1_strm0_data_valid  ;

  output                                          pe59__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane1_strm1_data_mask   ;
  input                                           std__pe59__lane1_strm1_data_valid  ;

  output                                          pe59__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane2_strm0_data_mask   ;
  input                                           std__pe59__lane2_strm0_data_valid  ;

  output                                          pe59__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane2_strm1_data_mask   ;
  input                                           std__pe59__lane2_strm1_data_valid  ;

  output                                          pe59__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane3_strm0_data_mask   ;
  input                                           std__pe59__lane3_strm0_data_valid  ;

  output                                          pe59__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane3_strm1_data_mask   ;
  input                                           std__pe59__lane3_strm1_data_valid  ;

  output                                          pe59__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane4_strm0_data_mask   ;
  input                                           std__pe59__lane4_strm0_data_valid  ;

  output                                          pe59__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane4_strm1_data_mask   ;
  input                                           std__pe59__lane4_strm1_data_valid  ;

  output                                          pe59__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane5_strm0_data_mask   ;
  input                                           std__pe59__lane5_strm0_data_valid  ;

  output                                          pe59__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane5_strm1_data_mask   ;
  input                                           std__pe59__lane5_strm1_data_valid  ;

  output                                          pe59__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane6_strm0_data_mask   ;
  input                                           std__pe59__lane6_strm0_data_valid  ;

  output                                          pe59__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane6_strm1_data_mask   ;
  input                                           std__pe59__lane6_strm1_data_valid  ;

  output                                          pe59__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane7_strm0_data_mask   ;
  input                                           std__pe59__lane7_strm0_data_valid  ;

  output                                          pe59__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane7_strm1_data_mask   ;
  input                                           std__pe59__lane7_strm1_data_valid  ;

  output                                          pe59__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane8_strm0_data_mask   ;
  input                                           std__pe59__lane8_strm0_data_valid  ;

  output                                          pe59__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane8_strm1_data_mask   ;
  input                                           std__pe59__lane8_strm1_data_valid  ;

  output                                          pe59__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane9_strm0_data_mask   ;
  input                                           std__pe59__lane9_strm0_data_valid  ;

  output                                          pe59__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane9_strm1_data_mask   ;
  input                                           std__pe59__lane9_strm1_data_valid  ;

  output                                          pe59__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane10_strm0_data_mask   ;
  input                                           std__pe59__lane10_strm0_data_valid  ;

  output                                          pe59__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane10_strm1_data_mask   ;
  input                                           std__pe59__lane10_strm1_data_valid  ;

  output                                          pe59__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane11_strm0_data_mask   ;
  input                                           std__pe59__lane11_strm0_data_valid  ;

  output                                          pe59__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane11_strm1_data_mask   ;
  input                                           std__pe59__lane11_strm1_data_valid  ;

  output                                          pe59__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane12_strm0_data_mask   ;
  input                                           std__pe59__lane12_strm0_data_valid  ;

  output                                          pe59__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane12_strm1_data_mask   ;
  input                                           std__pe59__lane12_strm1_data_valid  ;

  output                                          pe59__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane13_strm0_data_mask   ;
  input                                           std__pe59__lane13_strm0_data_valid  ;

  output                                          pe59__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane13_strm1_data_mask   ;
  input                                           std__pe59__lane13_strm1_data_valid  ;

  output                                          pe59__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane14_strm0_data_mask   ;
  input                                           std__pe59__lane14_strm0_data_valid  ;

  output                                          pe59__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane14_strm1_data_mask   ;
  input                                           std__pe59__lane14_strm1_data_valid  ;

  output                                          pe59__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane15_strm0_data_mask   ;
  input                                           std__pe59__lane15_strm0_data_valid  ;

  output                                          pe59__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane15_strm1_data_mask   ;
  input                                           std__pe59__lane15_strm1_data_valid  ;

  output                                          pe59__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane16_strm0_data_mask   ;
  input                                           std__pe59__lane16_strm0_data_valid  ;

  output                                          pe59__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane16_strm1_data_mask   ;
  input                                           std__pe59__lane16_strm1_data_valid  ;

  output                                          pe59__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane17_strm0_data_mask   ;
  input                                           std__pe59__lane17_strm0_data_valid  ;

  output                                          pe59__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane17_strm1_data_mask   ;
  input                                           std__pe59__lane17_strm1_data_valid  ;

  output                                          pe59__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane18_strm0_data_mask   ;
  input                                           std__pe59__lane18_strm0_data_valid  ;

  output                                          pe59__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane18_strm1_data_mask   ;
  input                                           std__pe59__lane18_strm1_data_valid  ;

  output                                          pe59__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane19_strm0_data_mask   ;
  input                                           std__pe59__lane19_strm0_data_valid  ;

  output                                          pe59__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane19_strm1_data_mask   ;
  input                                           std__pe59__lane19_strm1_data_valid  ;

  output                                          pe59__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane20_strm0_data_mask   ;
  input                                           std__pe59__lane20_strm0_data_valid  ;

  output                                          pe59__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane20_strm1_data_mask   ;
  input                                           std__pe59__lane20_strm1_data_valid  ;

  output                                          pe59__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane21_strm0_data_mask   ;
  input                                           std__pe59__lane21_strm0_data_valid  ;

  output                                          pe59__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane21_strm1_data_mask   ;
  input                                           std__pe59__lane21_strm1_data_valid  ;

  output                                          pe59__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane22_strm0_data_mask   ;
  input                                           std__pe59__lane22_strm0_data_valid  ;

  output                                          pe59__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane22_strm1_data_mask   ;
  input                                           std__pe59__lane22_strm1_data_valid  ;

  output                                          pe59__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane23_strm0_data_mask   ;
  input                                           std__pe59__lane23_strm0_data_valid  ;

  output                                          pe59__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane23_strm1_data_mask   ;
  input                                           std__pe59__lane23_strm1_data_valid  ;

  output                                          pe59__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane24_strm0_data_mask   ;
  input                                           std__pe59__lane24_strm0_data_valid  ;

  output                                          pe59__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane24_strm1_data_mask   ;
  input                                           std__pe59__lane24_strm1_data_valid  ;

  output                                          pe59__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane25_strm0_data_mask   ;
  input                                           std__pe59__lane25_strm0_data_valid  ;

  output                                          pe59__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane25_strm1_data_mask   ;
  input                                           std__pe59__lane25_strm1_data_valid  ;

  output                                          pe59__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane26_strm0_data_mask   ;
  input                                           std__pe59__lane26_strm0_data_valid  ;

  output                                          pe59__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane26_strm1_data_mask   ;
  input                                           std__pe59__lane26_strm1_data_valid  ;

  output                                          pe59__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane27_strm0_data_mask   ;
  input                                           std__pe59__lane27_strm0_data_valid  ;

  output                                          pe59__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane27_strm1_data_mask   ;
  input                                           std__pe59__lane27_strm1_data_valid  ;

  output                                          pe59__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane28_strm0_data_mask   ;
  input                                           std__pe59__lane28_strm0_data_valid  ;

  output                                          pe59__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane28_strm1_data_mask   ;
  input                                           std__pe59__lane28_strm1_data_valid  ;

  output                                          pe59__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane29_strm0_data_mask   ;
  input                                           std__pe59__lane29_strm0_data_valid  ;

  output                                          pe59__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane29_strm1_data_mask   ;
  input                                           std__pe59__lane29_strm1_data_valid  ;

  output                                          pe59__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane30_strm0_data_mask   ;
  input                                           std__pe59__lane30_strm0_data_valid  ;

  output                                          pe59__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane30_strm1_data_mask   ;
  input                                           std__pe59__lane30_strm1_data_valid  ;

  output                                          pe59__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane31_strm0_data_mask   ;
  input                                           std__pe59__lane31_strm0_data_valid  ;

  output                                          pe59__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe59__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe59__lane31_strm1_data_mask   ;
  input                                           std__pe59__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe60__peId                ;
  input                                         sys__pe60__allSynchronized     ;
  output                                        pe60__sys__thisSynchronized    ;
  output                                        pe60__sys__ready               ;
  output                                        pe60__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe60__oob_cntl            ;
  input                                         std__pe60__oob_valid           ;
  output                                        pe60__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe60__oob_type            ;
  output                                          pe60__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane0_strm0_data_mask   ;
  input                                           std__pe60__lane0_strm0_data_valid  ;

  output                                          pe60__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane0_strm1_data_mask   ;
  input                                           std__pe60__lane0_strm1_data_valid  ;

  output                                          pe60__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane1_strm0_data_mask   ;
  input                                           std__pe60__lane1_strm0_data_valid  ;

  output                                          pe60__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane1_strm1_data_mask   ;
  input                                           std__pe60__lane1_strm1_data_valid  ;

  output                                          pe60__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane2_strm0_data_mask   ;
  input                                           std__pe60__lane2_strm0_data_valid  ;

  output                                          pe60__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane2_strm1_data_mask   ;
  input                                           std__pe60__lane2_strm1_data_valid  ;

  output                                          pe60__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane3_strm0_data_mask   ;
  input                                           std__pe60__lane3_strm0_data_valid  ;

  output                                          pe60__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane3_strm1_data_mask   ;
  input                                           std__pe60__lane3_strm1_data_valid  ;

  output                                          pe60__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane4_strm0_data_mask   ;
  input                                           std__pe60__lane4_strm0_data_valid  ;

  output                                          pe60__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane4_strm1_data_mask   ;
  input                                           std__pe60__lane4_strm1_data_valid  ;

  output                                          pe60__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane5_strm0_data_mask   ;
  input                                           std__pe60__lane5_strm0_data_valid  ;

  output                                          pe60__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane5_strm1_data_mask   ;
  input                                           std__pe60__lane5_strm1_data_valid  ;

  output                                          pe60__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane6_strm0_data_mask   ;
  input                                           std__pe60__lane6_strm0_data_valid  ;

  output                                          pe60__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane6_strm1_data_mask   ;
  input                                           std__pe60__lane6_strm1_data_valid  ;

  output                                          pe60__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane7_strm0_data_mask   ;
  input                                           std__pe60__lane7_strm0_data_valid  ;

  output                                          pe60__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane7_strm1_data_mask   ;
  input                                           std__pe60__lane7_strm1_data_valid  ;

  output                                          pe60__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane8_strm0_data_mask   ;
  input                                           std__pe60__lane8_strm0_data_valid  ;

  output                                          pe60__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane8_strm1_data_mask   ;
  input                                           std__pe60__lane8_strm1_data_valid  ;

  output                                          pe60__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane9_strm0_data_mask   ;
  input                                           std__pe60__lane9_strm0_data_valid  ;

  output                                          pe60__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane9_strm1_data_mask   ;
  input                                           std__pe60__lane9_strm1_data_valid  ;

  output                                          pe60__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane10_strm0_data_mask   ;
  input                                           std__pe60__lane10_strm0_data_valid  ;

  output                                          pe60__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane10_strm1_data_mask   ;
  input                                           std__pe60__lane10_strm1_data_valid  ;

  output                                          pe60__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane11_strm0_data_mask   ;
  input                                           std__pe60__lane11_strm0_data_valid  ;

  output                                          pe60__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane11_strm1_data_mask   ;
  input                                           std__pe60__lane11_strm1_data_valid  ;

  output                                          pe60__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane12_strm0_data_mask   ;
  input                                           std__pe60__lane12_strm0_data_valid  ;

  output                                          pe60__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane12_strm1_data_mask   ;
  input                                           std__pe60__lane12_strm1_data_valid  ;

  output                                          pe60__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane13_strm0_data_mask   ;
  input                                           std__pe60__lane13_strm0_data_valid  ;

  output                                          pe60__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane13_strm1_data_mask   ;
  input                                           std__pe60__lane13_strm1_data_valid  ;

  output                                          pe60__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane14_strm0_data_mask   ;
  input                                           std__pe60__lane14_strm0_data_valid  ;

  output                                          pe60__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane14_strm1_data_mask   ;
  input                                           std__pe60__lane14_strm1_data_valid  ;

  output                                          pe60__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane15_strm0_data_mask   ;
  input                                           std__pe60__lane15_strm0_data_valid  ;

  output                                          pe60__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane15_strm1_data_mask   ;
  input                                           std__pe60__lane15_strm1_data_valid  ;

  output                                          pe60__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane16_strm0_data_mask   ;
  input                                           std__pe60__lane16_strm0_data_valid  ;

  output                                          pe60__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane16_strm1_data_mask   ;
  input                                           std__pe60__lane16_strm1_data_valid  ;

  output                                          pe60__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane17_strm0_data_mask   ;
  input                                           std__pe60__lane17_strm0_data_valid  ;

  output                                          pe60__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane17_strm1_data_mask   ;
  input                                           std__pe60__lane17_strm1_data_valid  ;

  output                                          pe60__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane18_strm0_data_mask   ;
  input                                           std__pe60__lane18_strm0_data_valid  ;

  output                                          pe60__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane18_strm1_data_mask   ;
  input                                           std__pe60__lane18_strm1_data_valid  ;

  output                                          pe60__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane19_strm0_data_mask   ;
  input                                           std__pe60__lane19_strm0_data_valid  ;

  output                                          pe60__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane19_strm1_data_mask   ;
  input                                           std__pe60__lane19_strm1_data_valid  ;

  output                                          pe60__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane20_strm0_data_mask   ;
  input                                           std__pe60__lane20_strm0_data_valid  ;

  output                                          pe60__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane20_strm1_data_mask   ;
  input                                           std__pe60__lane20_strm1_data_valid  ;

  output                                          pe60__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane21_strm0_data_mask   ;
  input                                           std__pe60__lane21_strm0_data_valid  ;

  output                                          pe60__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane21_strm1_data_mask   ;
  input                                           std__pe60__lane21_strm1_data_valid  ;

  output                                          pe60__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane22_strm0_data_mask   ;
  input                                           std__pe60__lane22_strm0_data_valid  ;

  output                                          pe60__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane22_strm1_data_mask   ;
  input                                           std__pe60__lane22_strm1_data_valid  ;

  output                                          pe60__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane23_strm0_data_mask   ;
  input                                           std__pe60__lane23_strm0_data_valid  ;

  output                                          pe60__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane23_strm1_data_mask   ;
  input                                           std__pe60__lane23_strm1_data_valid  ;

  output                                          pe60__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane24_strm0_data_mask   ;
  input                                           std__pe60__lane24_strm0_data_valid  ;

  output                                          pe60__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane24_strm1_data_mask   ;
  input                                           std__pe60__lane24_strm1_data_valid  ;

  output                                          pe60__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane25_strm0_data_mask   ;
  input                                           std__pe60__lane25_strm0_data_valid  ;

  output                                          pe60__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane25_strm1_data_mask   ;
  input                                           std__pe60__lane25_strm1_data_valid  ;

  output                                          pe60__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane26_strm0_data_mask   ;
  input                                           std__pe60__lane26_strm0_data_valid  ;

  output                                          pe60__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane26_strm1_data_mask   ;
  input                                           std__pe60__lane26_strm1_data_valid  ;

  output                                          pe60__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane27_strm0_data_mask   ;
  input                                           std__pe60__lane27_strm0_data_valid  ;

  output                                          pe60__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane27_strm1_data_mask   ;
  input                                           std__pe60__lane27_strm1_data_valid  ;

  output                                          pe60__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane28_strm0_data_mask   ;
  input                                           std__pe60__lane28_strm0_data_valid  ;

  output                                          pe60__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane28_strm1_data_mask   ;
  input                                           std__pe60__lane28_strm1_data_valid  ;

  output                                          pe60__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane29_strm0_data_mask   ;
  input                                           std__pe60__lane29_strm0_data_valid  ;

  output                                          pe60__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane29_strm1_data_mask   ;
  input                                           std__pe60__lane29_strm1_data_valid  ;

  output                                          pe60__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane30_strm0_data_mask   ;
  input                                           std__pe60__lane30_strm0_data_valid  ;

  output                                          pe60__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane30_strm1_data_mask   ;
  input                                           std__pe60__lane30_strm1_data_valid  ;

  output                                          pe60__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane31_strm0_data_mask   ;
  input                                           std__pe60__lane31_strm0_data_valid  ;

  output                                          pe60__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe60__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe60__lane31_strm1_data_mask   ;
  input                                           std__pe60__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe61__peId                ;
  input                                         sys__pe61__allSynchronized     ;
  output                                        pe61__sys__thisSynchronized    ;
  output                                        pe61__sys__ready               ;
  output                                        pe61__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe61__oob_cntl            ;
  input                                         std__pe61__oob_valid           ;
  output                                        pe61__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe61__oob_type            ;
  output                                          pe61__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane0_strm0_data_mask   ;
  input                                           std__pe61__lane0_strm0_data_valid  ;

  output                                          pe61__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane0_strm1_data_mask   ;
  input                                           std__pe61__lane0_strm1_data_valid  ;

  output                                          pe61__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane1_strm0_data_mask   ;
  input                                           std__pe61__lane1_strm0_data_valid  ;

  output                                          pe61__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane1_strm1_data_mask   ;
  input                                           std__pe61__lane1_strm1_data_valid  ;

  output                                          pe61__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane2_strm0_data_mask   ;
  input                                           std__pe61__lane2_strm0_data_valid  ;

  output                                          pe61__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane2_strm1_data_mask   ;
  input                                           std__pe61__lane2_strm1_data_valid  ;

  output                                          pe61__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane3_strm0_data_mask   ;
  input                                           std__pe61__lane3_strm0_data_valid  ;

  output                                          pe61__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane3_strm1_data_mask   ;
  input                                           std__pe61__lane3_strm1_data_valid  ;

  output                                          pe61__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane4_strm0_data_mask   ;
  input                                           std__pe61__lane4_strm0_data_valid  ;

  output                                          pe61__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane4_strm1_data_mask   ;
  input                                           std__pe61__lane4_strm1_data_valid  ;

  output                                          pe61__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane5_strm0_data_mask   ;
  input                                           std__pe61__lane5_strm0_data_valid  ;

  output                                          pe61__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane5_strm1_data_mask   ;
  input                                           std__pe61__lane5_strm1_data_valid  ;

  output                                          pe61__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane6_strm0_data_mask   ;
  input                                           std__pe61__lane6_strm0_data_valid  ;

  output                                          pe61__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane6_strm1_data_mask   ;
  input                                           std__pe61__lane6_strm1_data_valid  ;

  output                                          pe61__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane7_strm0_data_mask   ;
  input                                           std__pe61__lane7_strm0_data_valid  ;

  output                                          pe61__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane7_strm1_data_mask   ;
  input                                           std__pe61__lane7_strm1_data_valid  ;

  output                                          pe61__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane8_strm0_data_mask   ;
  input                                           std__pe61__lane8_strm0_data_valid  ;

  output                                          pe61__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane8_strm1_data_mask   ;
  input                                           std__pe61__lane8_strm1_data_valid  ;

  output                                          pe61__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane9_strm0_data_mask   ;
  input                                           std__pe61__lane9_strm0_data_valid  ;

  output                                          pe61__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane9_strm1_data_mask   ;
  input                                           std__pe61__lane9_strm1_data_valid  ;

  output                                          pe61__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane10_strm0_data_mask   ;
  input                                           std__pe61__lane10_strm0_data_valid  ;

  output                                          pe61__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane10_strm1_data_mask   ;
  input                                           std__pe61__lane10_strm1_data_valid  ;

  output                                          pe61__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane11_strm0_data_mask   ;
  input                                           std__pe61__lane11_strm0_data_valid  ;

  output                                          pe61__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane11_strm1_data_mask   ;
  input                                           std__pe61__lane11_strm1_data_valid  ;

  output                                          pe61__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane12_strm0_data_mask   ;
  input                                           std__pe61__lane12_strm0_data_valid  ;

  output                                          pe61__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane12_strm1_data_mask   ;
  input                                           std__pe61__lane12_strm1_data_valid  ;

  output                                          pe61__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane13_strm0_data_mask   ;
  input                                           std__pe61__lane13_strm0_data_valid  ;

  output                                          pe61__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane13_strm1_data_mask   ;
  input                                           std__pe61__lane13_strm1_data_valid  ;

  output                                          pe61__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane14_strm0_data_mask   ;
  input                                           std__pe61__lane14_strm0_data_valid  ;

  output                                          pe61__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane14_strm1_data_mask   ;
  input                                           std__pe61__lane14_strm1_data_valid  ;

  output                                          pe61__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane15_strm0_data_mask   ;
  input                                           std__pe61__lane15_strm0_data_valid  ;

  output                                          pe61__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane15_strm1_data_mask   ;
  input                                           std__pe61__lane15_strm1_data_valid  ;

  output                                          pe61__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane16_strm0_data_mask   ;
  input                                           std__pe61__lane16_strm0_data_valid  ;

  output                                          pe61__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane16_strm1_data_mask   ;
  input                                           std__pe61__lane16_strm1_data_valid  ;

  output                                          pe61__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane17_strm0_data_mask   ;
  input                                           std__pe61__lane17_strm0_data_valid  ;

  output                                          pe61__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane17_strm1_data_mask   ;
  input                                           std__pe61__lane17_strm1_data_valid  ;

  output                                          pe61__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane18_strm0_data_mask   ;
  input                                           std__pe61__lane18_strm0_data_valid  ;

  output                                          pe61__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane18_strm1_data_mask   ;
  input                                           std__pe61__lane18_strm1_data_valid  ;

  output                                          pe61__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane19_strm0_data_mask   ;
  input                                           std__pe61__lane19_strm0_data_valid  ;

  output                                          pe61__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane19_strm1_data_mask   ;
  input                                           std__pe61__lane19_strm1_data_valid  ;

  output                                          pe61__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane20_strm0_data_mask   ;
  input                                           std__pe61__lane20_strm0_data_valid  ;

  output                                          pe61__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane20_strm1_data_mask   ;
  input                                           std__pe61__lane20_strm1_data_valid  ;

  output                                          pe61__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane21_strm0_data_mask   ;
  input                                           std__pe61__lane21_strm0_data_valid  ;

  output                                          pe61__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane21_strm1_data_mask   ;
  input                                           std__pe61__lane21_strm1_data_valid  ;

  output                                          pe61__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane22_strm0_data_mask   ;
  input                                           std__pe61__lane22_strm0_data_valid  ;

  output                                          pe61__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane22_strm1_data_mask   ;
  input                                           std__pe61__lane22_strm1_data_valid  ;

  output                                          pe61__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane23_strm0_data_mask   ;
  input                                           std__pe61__lane23_strm0_data_valid  ;

  output                                          pe61__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane23_strm1_data_mask   ;
  input                                           std__pe61__lane23_strm1_data_valid  ;

  output                                          pe61__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane24_strm0_data_mask   ;
  input                                           std__pe61__lane24_strm0_data_valid  ;

  output                                          pe61__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane24_strm1_data_mask   ;
  input                                           std__pe61__lane24_strm1_data_valid  ;

  output                                          pe61__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane25_strm0_data_mask   ;
  input                                           std__pe61__lane25_strm0_data_valid  ;

  output                                          pe61__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane25_strm1_data_mask   ;
  input                                           std__pe61__lane25_strm1_data_valid  ;

  output                                          pe61__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane26_strm0_data_mask   ;
  input                                           std__pe61__lane26_strm0_data_valid  ;

  output                                          pe61__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane26_strm1_data_mask   ;
  input                                           std__pe61__lane26_strm1_data_valid  ;

  output                                          pe61__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane27_strm0_data_mask   ;
  input                                           std__pe61__lane27_strm0_data_valid  ;

  output                                          pe61__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane27_strm1_data_mask   ;
  input                                           std__pe61__lane27_strm1_data_valid  ;

  output                                          pe61__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane28_strm0_data_mask   ;
  input                                           std__pe61__lane28_strm0_data_valid  ;

  output                                          pe61__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane28_strm1_data_mask   ;
  input                                           std__pe61__lane28_strm1_data_valid  ;

  output                                          pe61__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane29_strm0_data_mask   ;
  input                                           std__pe61__lane29_strm0_data_valid  ;

  output                                          pe61__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane29_strm1_data_mask   ;
  input                                           std__pe61__lane29_strm1_data_valid  ;

  output                                          pe61__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane30_strm0_data_mask   ;
  input                                           std__pe61__lane30_strm0_data_valid  ;

  output                                          pe61__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane30_strm1_data_mask   ;
  input                                           std__pe61__lane30_strm1_data_valid  ;

  output                                          pe61__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane31_strm0_data_mask   ;
  input                                           std__pe61__lane31_strm0_data_valid  ;

  output                                          pe61__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe61__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe61__lane31_strm1_data_mask   ;
  input                                           std__pe61__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe62__peId                ;
  input                                         sys__pe62__allSynchronized     ;
  output                                        pe62__sys__thisSynchronized    ;
  output                                        pe62__sys__ready               ;
  output                                        pe62__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe62__oob_cntl            ;
  input                                         std__pe62__oob_valid           ;
  output                                        pe62__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe62__oob_type            ;
  output                                          pe62__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane0_strm0_data_mask   ;
  input                                           std__pe62__lane0_strm0_data_valid  ;

  output                                          pe62__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane0_strm1_data_mask   ;
  input                                           std__pe62__lane0_strm1_data_valid  ;

  output                                          pe62__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane1_strm0_data_mask   ;
  input                                           std__pe62__lane1_strm0_data_valid  ;

  output                                          pe62__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane1_strm1_data_mask   ;
  input                                           std__pe62__lane1_strm1_data_valid  ;

  output                                          pe62__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane2_strm0_data_mask   ;
  input                                           std__pe62__lane2_strm0_data_valid  ;

  output                                          pe62__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane2_strm1_data_mask   ;
  input                                           std__pe62__lane2_strm1_data_valid  ;

  output                                          pe62__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane3_strm0_data_mask   ;
  input                                           std__pe62__lane3_strm0_data_valid  ;

  output                                          pe62__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane3_strm1_data_mask   ;
  input                                           std__pe62__lane3_strm1_data_valid  ;

  output                                          pe62__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane4_strm0_data_mask   ;
  input                                           std__pe62__lane4_strm0_data_valid  ;

  output                                          pe62__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane4_strm1_data_mask   ;
  input                                           std__pe62__lane4_strm1_data_valid  ;

  output                                          pe62__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane5_strm0_data_mask   ;
  input                                           std__pe62__lane5_strm0_data_valid  ;

  output                                          pe62__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane5_strm1_data_mask   ;
  input                                           std__pe62__lane5_strm1_data_valid  ;

  output                                          pe62__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane6_strm0_data_mask   ;
  input                                           std__pe62__lane6_strm0_data_valid  ;

  output                                          pe62__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane6_strm1_data_mask   ;
  input                                           std__pe62__lane6_strm1_data_valid  ;

  output                                          pe62__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane7_strm0_data_mask   ;
  input                                           std__pe62__lane7_strm0_data_valid  ;

  output                                          pe62__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane7_strm1_data_mask   ;
  input                                           std__pe62__lane7_strm1_data_valid  ;

  output                                          pe62__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane8_strm0_data_mask   ;
  input                                           std__pe62__lane8_strm0_data_valid  ;

  output                                          pe62__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane8_strm1_data_mask   ;
  input                                           std__pe62__lane8_strm1_data_valid  ;

  output                                          pe62__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane9_strm0_data_mask   ;
  input                                           std__pe62__lane9_strm0_data_valid  ;

  output                                          pe62__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane9_strm1_data_mask   ;
  input                                           std__pe62__lane9_strm1_data_valid  ;

  output                                          pe62__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane10_strm0_data_mask   ;
  input                                           std__pe62__lane10_strm0_data_valid  ;

  output                                          pe62__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane10_strm1_data_mask   ;
  input                                           std__pe62__lane10_strm1_data_valid  ;

  output                                          pe62__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane11_strm0_data_mask   ;
  input                                           std__pe62__lane11_strm0_data_valid  ;

  output                                          pe62__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane11_strm1_data_mask   ;
  input                                           std__pe62__lane11_strm1_data_valid  ;

  output                                          pe62__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane12_strm0_data_mask   ;
  input                                           std__pe62__lane12_strm0_data_valid  ;

  output                                          pe62__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane12_strm1_data_mask   ;
  input                                           std__pe62__lane12_strm1_data_valid  ;

  output                                          pe62__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane13_strm0_data_mask   ;
  input                                           std__pe62__lane13_strm0_data_valid  ;

  output                                          pe62__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane13_strm1_data_mask   ;
  input                                           std__pe62__lane13_strm1_data_valid  ;

  output                                          pe62__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane14_strm0_data_mask   ;
  input                                           std__pe62__lane14_strm0_data_valid  ;

  output                                          pe62__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane14_strm1_data_mask   ;
  input                                           std__pe62__lane14_strm1_data_valid  ;

  output                                          pe62__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane15_strm0_data_mask   ;
  input                                           std__pe62__lane15_strm0_data_valid  ;

  output                                          pe62__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane15_strm1_data_mask   ;
  input                                           std__pe62__lane15_strm1_data_valid  ;

  output                                          pe62__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane16_strm0_data_mask   ;
  input                                           std__pe62__lane16_strm0_data_valid  ;

  output                                          pe62__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane16_strm1_data_mask   ;
  input                                           std__pe62__lane16_strm1_data_valid  ;

  output                                          pe62__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane17_strm0_data_mask   ;
  input                                           std__pe62__lane17_strm0_data_valid  ;

  output                                          pe62__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane17_strm1_data_mask   ;
  input                                           std__pe62__lane17_strm1_data_valid  ;

  output                                          pe62__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane18_strm0_data_mask   ;
  input                                           std__pe62__lane18_strm0_data_valid  ;

  output                                          pe62__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane18_strm1_data_mask   ;
  input                                           std__pe62__lane18_strm1_data_valid  ;

  output                                          pe62__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane19_strm0_data_mask   ;
  input                                           std__pe62__lane19_strm0_data_valid  ;

  output                                          pe62__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane19_strm1_data_mask   ;
  input                                           std__pe62__lane19_strm1_data_valid  ;

  output                                          pe62__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane20_strm0_data_mask   ;
  input                                           std__pe62__lane20_strm0_data_valid  ;

  output                                          pe62__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane20_strm1_data_mask   ;
  input                                           std__pe62__lane20_strm1_data_valid  ;

  output                                          pe62__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane21_strm0_data_mask   ;
  input                                           std__pe62__lane21_strm0_data_valid  ;

  output                                          pe62__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane21_strm1_data_mask   ;
  input                                           std__pe62__lane21_strm1_data_valid  ;

  output                                          pe62__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane22_strm0_data_mask   ;
  input                                           std__pe62__lane22_strm0_data_valid  ;

  output                                          pe62__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane22_strm1_data_mask   ;
  input                                           std__pe62__lane22_strm1_data_valid  ;

  output                                          pe62__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane23_strm0_data_mask   ;
  input                                           std__pe62__lane23_strm0_data_valid  ;

  output                                          pe62__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane23_strm1_data_mask   ;
  input                                           std__pe62__lane23_strm1_data_valid  ;

  output                                          pe62__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane24_strm0_data_mask   ;
  input                                           std__pe62__lane24_strm0_data_valid  ;

  output                                          pe62__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane24_strm1_data_mask   ;
  input                                           std__pe62__lane24_strm1_data_valid  ;

  output                                          pe62__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane25_strm0_data_mask   ;
  input                                           std__pe62__lane25_strm0_data_valid  ;

  output                                          pe62__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane25_strm1_data_mask   ;
  input                                           std__pe62__lane25_strm1_data_valid  ;

  output                                          pe62__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane26_strm0_data_mask   ;
  input                                           std__pe62__lane26_strm0_data_valid  ;

  output                                          pe62__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane26_strm1_data_mask   ;
  input                                           std__pe62__lane26_strm1_data_valid  ;

  output                                          pe62__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane27_strm0_data_mask   ;
  input                                           std__pe62__lane27_strm0_data_valid  ;

  output                                          pe62__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane27_strm1_data_mask   ;
  input                                           std__pe62__lane27_strm1_data_valid  ;

  output                                          pe62__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane28_strm0_data_mask   ;
  input                                           std__pe62__lane28_strm0_data_valid  ;

  output                                          pe62__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane28_strm1_data_mask   ;
  input                                           std__pe62__lane28_strm1_data_valid  ;

  output                                          pe62__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane29_strm0_data_mask   ;
  input                                           std__pe62__lane29_strm0_data_valid  ;

  output                                          pe62__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane29_strm1_data_mask   ;
  input                                           std__pe62__lane29_strm1_data_valid  ;

  output                                          pe62__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane30_strm0_data_mask   ;
  input                                           std__pe62__lane30_strm0_data_valid  ;

  output                                          pe62__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane30_strm1_data_mask   ;
  input                                           std__pe62__lane30_strm1_data_valid  ;

  output                                          pe62__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane31_strm0_data_mask   ;
  input                                           std__pe62__lane31_strm0_data_valid  ;

  output                                          pe62__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe62__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe62__lane31_strm1_data_mask   ;
  input                                           std__pe62__lane31_strm1_data_valid  ;

  // General control and status                                                  
  input [`PE_PE_ID_RANGE                 ]      sys__pe63__peId                ;
  input                                         sys__pe63__allSynchronized     ;
  output                                        pe63__sys__thisSynchronized    ;
  output                                        pe63__sys__ready               ;
  output                                        pe63__sys__complete            ;
  // OOB controls how the lanes are interpreted                                  
  input [`COMMON_STD_INTF_CNTL_RANGE     ]      std__pe63__oob_cntl            ;
  input                                         std__pe63__oob_valid           ;
  output                                        pe63__std__oob_ready           ;
  input [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      std__pe63__oob_type            ;
  output                                          pe63__std__lane0_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane0_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane0_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane0_strm0_data_mask   ;
  input                                           std__pe63__lane0_strm0_data_valid  ;

  output                                          pe63__std__lane0_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane0_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane0_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane0_strm1_data_mask   ;
  input                                           std__pe63__lane0_strm1_data_valid  ;

  output                                          pe63__std__lane1_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane1_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane1_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane1_strm0_data_mask   ;
  input                                           std__pe63__lane1_strm0_data_valid  ;

  output                                          pe63__std__lane1_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane1_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane1_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane1_strm1_data_mask   ;
  input                                           std__pe63__lane1_strm1_data_valid  ;

  output                                          pe63__std__lane2_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane2_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane2_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane2_strm0_data_mask   ;
  input                                           std__pe63__lane2_strm0_data_valid  ;

  output                                          pe63__std__lane2_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane2_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane2_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane2_strm1_data_mask   ;
  input                                           std__pe63__lane2_strm1_data_valid  ;

  output                                          pe63__std__lane3_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane3_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane3_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane3_strm0_data_mask   ;
  input                                           std__pe63__lane3_strm0_data_valid  ;

  output                                          pe63__std__lane3_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane3_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane3_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane3_strm1_data_mask   ;
  input                                           std__pe63__lane3_strm1_data_valid  ;

  output                                          pe63__std__lane4_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane4_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane4_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane4_strm0_data_mask   ;
  input                                           std__pe63__lane4_strm0_data_valid  ;

  output                                          pe63__std__lane4_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane4_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane4_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane4_strm1_data_mask   ;
  input                                           std__pe63__lane4_strm1_data_valid  ;

  output                                          pe63__std__lane5_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane5_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane5_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane5_strm0_data_mask   ;
  input                                           std__pe63__lane5_strm0_data_valid  ;

  output                                          pe63__std__lane5_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane5_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane5_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane5_strm1_data_mask   ;
  input                                           std__pe63__lane5_strm1_data_valid  ;

  output                                          pe63__std__lane6_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane6_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane6_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane6_strm0_data_mask   ;
  input                                           std__pe63__lane6_strm0_data_valid  ;

  output                                          pe63__std__lane6_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane6_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane6_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane6_strm1_data_mask   ;
  input                                           std__pe63__lane6_strm1_data_valid  ;

  output                                          pe63__std__lane7_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane7_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane7_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane7_strm0_data_mask   ;
  input                                           std__pe63__lane7_strm0_data_valid  ;

  output                                          pe63__std__lane7_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane7_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane7_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane7_strm1_data_mask   ;
  input                                           std__pe63__lane7_strm1_data_valid  ;

  output                                          pe63__std__lane8_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane8_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane8_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane8_strm0_data_mask   ;
  input                                           std__pe63__lane8_strm0_data_valid  ;

  output                                          pe63__std__lane8_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane8_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane8_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane8_strm1_data_mask   ;
  input                                           std__pe63__lane8_strm1_data_valid  ;

  output                                          pe63__std__lane9_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane9_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane9_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane9_strm0_data_mask   ;
  input                                           std__pe63__lane9_strm0_data_valid  ;

  output                                          pe63__std__lane9_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane9_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane9_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane9_strm1_data_mask   ;
  input                                           std__pe63__lane9_strm1_data_valid  ;

  output                                          pe63__std__lane10_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane10_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane10_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane10_strm0_data_mask   ;
  input                                           std__pe63__lane10_strm0_data_valid  ;

  output                                          pe63__std__lane10_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane10_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane10_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane10_strm1_data_mask   ;
  input                                           std__pe63__lane10_strm1_data_valid  ;

  output                                          pe63__std__lane11_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane11_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane11_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane11_strm0_data_mask   ;
  input                                           std__pe63__lane11_strm0_data_valid  ;

  output                                          pe63__std__lane11_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane11_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane11_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane11_strm1_data_mask   ;
  input                                           std__pe63__lane11_strm1_data_valid  ;

  output                                          pe63__std__lane12_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane12_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane12_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane12_strm0_data_mask   ;
  input                                           std__pe63__lane12_strm0_data_valid  ;

  output                                          pe63__std__lane12_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane12_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane12_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane12_strm1_data_mask   ;
  input                                           std__pe63__lane12_strm1_data_valid  ;

  output                                          pe63__std__lane13_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane13_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane13_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane13_strm0_data_mask   ;
  input                                           std__pe63__lane13_strm0_data_valid  ;

  output                                          pe63__std__lane13_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane13_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane13_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane13_strm1_data_mask   ;
  input                                           std__pe63__lane13_strm1_data_valid  ;

  output                                          pe63__std__lane14_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane14_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane14_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane14_strm0_data_mask   ;
  input                                           std__pe63__lane14_strm0_data_valid  ;

  output                                          pe63__std__lane14_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane14_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane14_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane14_strm1_data_mask   ;
  input                                           std__pe63__lane14_strm1_data_valid  ;

  output                                          pe63__std__lane15_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane15_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane15_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane15_strm0_data_mask   ;
  input                                           std__pe63__lane15_strm0_data_valid  ;

  output                                          pe63__std__lane15_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane15_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane15_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane15_strm1_data_mask   ;
  input                                           std__pe63__lane15_strm1_data_valid  ;

  output                                          pe63__std__lane16_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane16_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane16_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane16_strm0_data_mask   ;
  input                                           std__pe63__lane16_strm0_data_valid  ;

  output                                          pe63__std__lane16_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane16_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane16_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane16_strm1_data_mask   ;
  input                                           std__pe63__lane16_strm1_data_valid  ;

  output                                          pe63__std__lane17_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane17_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane17_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane17_strm0_data_mask   ;
  input                                           std__pe63__lane17_strm0_data_valid  ;

  output                                          pe63__std__lane17_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane17_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane17_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane17_strm1_data_mask   ;
  input                                           std__pe63__lane17_strm1_data_valid  ;

  output                                          pe63__std__lane18_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane18_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane18_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane18_strm0_data_mask   ;
  input                                           std__pe63__lane18_strm0_data_valid  ;

  output                                          pe63__std__lane18_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane18_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane18_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane18_strm1_data_mask   ;
  input                                           std__pe63__lane18_strm1_data_valid  ;

  output                                          pe63__std__lane19_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane19_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane19_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane19_strm0_data_mask   ;
  input                                           std__pe63__lane19_strm0_data_valid  ;

  output                                          pe63__std__lane19_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane19_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane19_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane19_strm1_data_mask   ;
  input                                           std__pe63__lane19_strm1_data_valid  ;

  output                                          pe63__std__lane20_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane20_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane20_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane20_strm0_data_mask   ;
  input                                           std__pe63__lane20_strm0_data_valid  ;

  output                                          pe63__std__lane20_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane20_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane20_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane20_strm1_data_mask   ;
  input                                           std__pe63__lane20_strm1_data_valid  ;

  output                                          pe63__std__lane21_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane21_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane21_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane21_strm0_data_mask   ;
  input                                           std__pe63__lane21_strm0_data_valid  ;

  output                                          pe63__std__lane21_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane21_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane21_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane21_strm1_data_mask   ;
  input                                           std__pe63__lane21_strm1_data_valid  ;

  output                                          pe63__std__lane22_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane22_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane22_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane22_strm0_data_mask   ;
  input                                           std__pe63__lane22_strm0_data_valid  ;

  output                                          pe63__std__lane22_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane22_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane22_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane22_strm1_data_mask   ;
  input                                           std__pe63__lane22_strm1_data_valid  ;

  output                                          pe63__std__lane23_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane23_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane23_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane23_strm0_data_mask   ;
  input                                           std__pe63__lane23_strm0_data_valid  ;

  output                                          pe63__std__lane23_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane23_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane23_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane23_strm1_data_mask   ;
  input                                           std__pe63__lane23_strm1_data_valid  ;

  output                                          pe63__std__lane24_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane24_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane24_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane24_strm0_data_mask   ;
  input                                           std__pe63__lane24_strm0_data_valid  ;

  output                                          pe63__std__lane24_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane24_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane24_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane24_strm1_data_mask   ;
  input                                           std__pe63__lane24_strm1_data_valid  ;

  output                                          pe63__std__lane25_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane25_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane25_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane25_strm0_data_mask   ;
  input                                           std__pe63__lane25_strm0_data_valid  ;

  output                                          pe63__std__lane25_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane25_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane25_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane25_strm1_data_mask   ;
  input                                           std__pe63__lane25_strm1_data_valid  ;

  output                                          pe63__std__lane26_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane26_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane26_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane26_strm0_data_mask   ;
  input                                           std__pe63__lane26_strm0_data_valid  ;

  output                                          pe63__std__lane26_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane26_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane26_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane26_strm1_data_mask   ;
  input                                           std__pe63__lane26_strm1_data_valid  ;

  output                                          pe63__std__lane27_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane27_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane27_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane27_strm0_data_mask   ;
  input                                           std__pe63__lane27_strm0_data_valid  ;

  output                                          pe63__std__lane27_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane27_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane27_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane27_strm1_data_mask   ;
  input                                           std__pe63__lane27_strm1_data_valid  ;

  output                                          pe63__std__lane28_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane28_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane28_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane28_strm0_data_mask   ;
  input                                           std__pe63__lane28_strm0_data_valid  ;

  output                                          pe63__std__lane28_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane28_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane28_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane28_strm1_data_mask   ;
  input                                           std__pe63__lane28_strm1_data_valid  ;

  output                                          pe63__std__lane29_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane29_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane29_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane29_strm0_data_mask   ;
  input                                           std__pe63__lane29_strm0_data_valid  ;

  output                                          pe63__std__lane29_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane29_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane29_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane29_strm1_data_mask   ;
  input                                           std__pe63__lane29_strm1_data_valid  ;

  output                                          pe63__std__lane30_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane30_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane30_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane30_strm0_data_mask   ;
  input                                           std__pe63__lane30_strm0_data_valid  ;

  output                                          pe63__std__lane30_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane30_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane30_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane30_strm1_data_mask   ;
  input                                           std__pe63__lane30_strm1_data_valid  ;

  output                                          pe63__std__lane31_strm0_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane31_strm0_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane31_strm0_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane31_strm0_data_mask   ;
  input                                           std__pe63__lane31_strm0_data_valid  ;

  output                                          pe63__std__lane31_strm1_ready       ;
  input [`COMMON_STD_INTF_CNTL_RANGE      ]       std__pe63__lane31_strm1_cntl        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane31_strm1_data        ;
  input [`STACK_DOWN_INTF_STRM_DATA_RANGE ]       std__pe63__lane31_strm1_data_mask   ;
  input                                           std__pe63__lane31_strm1_data_valid  ;
