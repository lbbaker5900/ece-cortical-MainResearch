
            .stu__mgr0__valid        ( stu__mgr0__valid     ),
            .stu__mgr0__cntl         ( stu__mgr0__cntl      ),
            .mgr0__stu__ready        ( mgr0__stu__ready     ),
            .stu__mgr0__type         ( stu__mgr0__type      ),
            .stu__mgr0__data         ( stu__mgr0__data      ),
            .stu__mgr0__oob_data     ( stu__mgr0__oob_data  ),

            .stu__mgr1__valid        ( stu__mgr1__valid     ),
            .stu__mgr1__cntl         ( stu__mgr1__cntl      ),
            .mgr1__stu__ready        ( mgr1__stu__ready     ),
            .stu__mgr1__type         ( stu__mgr1__type      ),
            .stu__mgr1__data         ( stu__mgr1__data      ),
            .stu__mgr1__oob_data     ( stu__mgr1__oob_data  ),

            .stu__mgr2__valid        ( stu__mgr2__valid     ),
            .stu__mgr2__cntl         ( stu__mgr2__cntl      ),
            .mgr2__stu__ready        ( mgr2__stu__ready     ),
            .stu__mgr2__type         ( stu__mgr2__type      ),
            .stu__mgr2__data         ( stu__mgr2__data      ),
            .stu__mgr2__oob_data     ( stu__mgr2__oob_data  ),

            .stu__mgr3__valid        ( stu__mgr3__valid     ),
            .stu__mgr3__cntl         ( stu__mgr3__cntl      ),
            .mgr3__stu__ready        ( mgr3__stu__ready     ),
            .stu__mgr3__type         ( stu__mgr3__type      ),
            .stu__mgr3__data         ( stu__mgr3__data      ),
            .stu__mgr3__oob_data     ( stu__mgr3__oob_data  ),

            .stu__mgr4__valid        ( stu__mgr4__valid     ),
            .stu__mgr4__cntl         ( stu__mgr4__cntl      ),
            .mgr4__stu__ready        ( mgr4__stu__ready     ),
            .stu__mgr4__type         ( stu__mgr4__type      ),
            .stu__mgr4__data         ( stu__mgr4__data      ),
            .stu__mgr4__oob_data     ( stu__mgr4__oob_data  ),

            .stu__mgr5__valid        ( stu__mgr5__valid     ),
            .stu__mgr5__cntl         ( stu__mgr5__cntl      ),
            .mgr5__stu__ready        ( mgr5__stu__ready     ),
            .stu__mgr5__type         ( stu__mgr5__type      ),
            .stu__mgr5__data         ( stu__mgr5__data      ),
            .stu__mgr5__oob_data     ( stu__mgr5__oob_data  ),

            .stu__mgr6__valid        ( stu__mgr6__valid     ),
            .stu__mgr6__cntl         ( stu__mgr6__cntl      ),
            .mgr6__stu__ready        ( mgr6__stu__ready     ),
            .stu__mgr6__type         ( stu__mgr6__type      ),
            .stu__mgr6__data         ( stu__mgr6__data      ),
            .stu__mgr6__oob_data     ( stu__mgr6__oob_data  ),

            .stu__mgr7__valid        ( stu__mgr7__valid     ),
            .stu__mgr7__cntl         ( stu__mgr7__cntl      ),
            .mgr7__stu__ready        ( mgr7__stu__ready     ),
            .stu__mgr7__type         ( stu__mgr7__type      ),
            .stu__mgr7__data         ( stu__mgr7__data      ),
            .stu__mgr7__oob_data     ( stu__mgr7__oob_data  ),

            .stu__mgr8__valid        ( stu__mgr8__valid     ),
            .stu__mgr8__cntl         ( stu__mgr8__cntl      ),
            .mgr8__stu__ready        ( mgr8__stu__ready     ),
            .stu__mgr8__type         ( stu__mgr8__type      ),
            .stu__mgr8__data         ( stu__mgr8__data      ),
            .stu__mgr8__oob_data     ( stu__mgr8__oob_data  ),

            .stu__mgr9__valid        ( stu__mgr9__valid     ),
            .stu__mgr9__cntl         ( stu__mgr9__cntl      ),
            .mgr9__stu__ready        ( mgr9__stu__ready     ),
            .stu__mgr9__type         ( stu__mgr9__type      ),
            .stu__mgr9__data         ( stu__mgr9__data      ),
            .stu__mgr9__oob_data     ( stu__mgr9__oob_data  ),

            .stu__mgr10__valid        ( stu__mgr10__valid     ),
            .stu__mgr10__cntl         ( stu__mgr10__cntl      ),
            .mgr10__stu__ready        ( mgr10__stu__ready     ),
            .stu__mgr10__type         ( stu__mgr10__type      ),
            .stu__mgr10__data         ( stu__mgr10__data      ),
            .stu__mgr10__oob_data     ( stu__mgr10__oob_data  ),

            .stu__mgr11__valid        ( stu__mgr11__valid     ),
            .stu__mgr11__cntl         ( stu__mgr11__cntl      ),
            .mgr11__stu__ready        ( mgr11__stu__ready     ),
            .stu__mgr11__type         ( stu__mgr11__type      ),
            .stu__mgr11__data         ( stu__mgr11__data      ),
            .stu__mgr11__oob_data     ( stu__mgr11__oob_data  ),

            .stu__mgr12__valid        ( stu__mgr12__valid     ),
            .stu__mgr12__cntl         ( stu__mgr12__cntl      ),
            .mgr12__stu__ready        ( mgr12__stu__ready     ),
            .stu__mgr12__type         ( stu__mgr12__type      ),
            .stu__mgr12__data         ( stu__mgr12__data      ),
            .stu__mgr12__oob_data     ( stu__mgr12__oob_data  ),

            .stu__mgr13__valid        ( stu__mgr13__valid     ),
            .stu__mgr13__cntl         ( stu__mgr13__cntl      ),
            .mgr13__stu__ready        ( mgr13__stu__ready     ),
            .stu__mgr13__type         ( stu__mgr13__type      ),
            .stu__mgr13__data         ( stu__mgr13__data      ),
            .stu__mgr13__oob_data     ( stu__mgr13__oob_data  ),

            .stu__mgr14__valid        ( stu__mgr14__valid     ),
            .stu__mgr14__cntl         ( stu__mgr14__cntl      ),
            .mgr14__stu__ready        ( mgr14__stu__ready     ),
            .stu__mgr14__type         ( stu__mgr14__type      ),
            .stu__mgr14__data         ( stu__mgr14__data      ),
            .stu__mgr14__oob_data     ( stu__mgr14__oob_data  ),

            .stu__mgr15__valid        ( stu__mgr15__valid     ),
            .stu__mgr15__cntl         ( stu__mgr15__cntl      ),
            .mgr15__stu__ready        ( mgr15__stu__ready     ),
            .stu__mgr15__type         ( stu__mgr15__type      ),
            .stu__mgr15__data         ( stu__mgr15__data      ),
            .stu__mgr15__oob_data     ( stu__mgr15__oob_data  ),

            .stu__mgr16__valid        ( stu__mgr16__valid     ),
            .stu__mgr16__cntl         ( stu__mgr16__cntl      ),
            .mgr16__stu__ready        ( mgr16__stu__ready     ),
            .stu__mgr16__type         ( stu__mgr16__type      ),
            .stu__mgr16__data         ( stu__mgr16__data      ),
            .stu__mgr16__oob_data     ( stu__mgr16__oob_data  ),

            .stu__mgr17__valid        ( stu__mgr17__valid     ),
            .stu__mgr17__cntl         ( stu__mgr17__cntl      ),
            .mgr17__stu__ready        ( mgr17__stu__ready     ),
            .stu__mgr17__type         ( stu__mgr17__type      ),
            .stu__mgr17__data         ( stu__mgr17__data      ),
            .stu__mgr17__oob_data     ( stu__mgr17__oob_data  ),

            .stu__mgr18__valid        ( stu__mgr18__valid     ),
            .stu__mgr18__cntl         ( stu__mgr18__cntl      ),
            .mgr18__stu__ready        ( mgr18__stu__ready     ),
            .stu__mgr18__type         ( stu__mgr18__type      ),
            .stu__mgr18__data         ( stu__mgr18__data      ),
            .stu__mgr18__oob_data     ( stu__mgr18__oob_data  ),

            .stu__mgr19__valid        ( stu__mgr19__valid     ),
            .stu__mgr19__cntl         ( stu__mgr19__cntl      ),
            .mgr19__stu__ready        ( mgr19__stu__ready     ),
            .stu__mgr19__type         ( stu__mgr19__type      ),
            .stu__mgr19__data         ( stu__mgr19__data      ),
            .stu__mgr19__oob_data     ( stu__mgr19__oob_data  ),

            .stu__mgr20__valid        ( stu__mgr20__valid     ),
            .stu__mgr20__cntl         ( stu__mgr20__cntl      ),
            .mgr20__stu__ready        ( mgr20__stu__ready     ),
            .stu__mgr20__type         ( stu__mgr20__type      ),
            .stu__mgr20__data         ( stu__mgr20__data      ),
            .stu__mgr20__oob_data     ( stu__mgr20__oob_data  ),

            .stu__mgr21__valid        ( stu__mgr21__valid     ),
            .stu__mgr21__cntl         ( stu__mgr21__cntl      ),
            .mgr21__stu__ready        ( mgr21__stu__ready     ),
            .stu__mgr21__type         ( stu__mgr21__type      ),
            .stu__mgr21__data         ( stu__mgr21__data      ),
            .stu__mgr21__oob_data     ( stu__mgr21__oob_data  ),

            .stu__mgr22__valid        ( stu__mgr22__valid     ),
            .stu__mgr22__cntl         ( stu__mgr22__cntl      ),
            .mgr22__stu__ready        ( mgr22__stu__ready     ),
            .stu__mgr22__type         ( stu__mgr22__type      ),
            .stu__mgr22__data         ( stu__mgr22__data      ),
            .stu__mgr22__oob_data     ( stu__mgr22__oob_data  ),

            .stu__mgr23__valid        ( stu__mgr23__valid     ),
            .stu__mgr23__cntl         ( stu__mgr23__cntl      ),
            .mgr23__stu__ready        ( mgr23__stu__ready     ),
            .stu__mgr23__type         ( stu__mgr23__type      ),
            .stu__mgr23__data         ( stu__mgr23__data      ),
            .stu__mgr23__oob_data     ( stu__mgr23__oob_data  ),

            .stu__mgr24__valid        ( stu__mgr24__valid     ),
            .stu__mgr24__cntl         ( stu__mgr24__cntl      ),
            .mgr24__stu__ready        ( mgr24__stu__ready     ),
            .stu__mgr24__type         ( stu__mgr24__type      ),
            .stu__mgr24__data         ( stu__mgr24__data      ),
            .stu__mgr24__oob_data     ( stu__mgr24__oob_data  ),

            .stu__mgr25__valid        ( stu__mgr25__valid     ),
            .stu__mgr25__cntl         ( stu__mgr25__cntl      ),
            .mgr25__stu__ready        ( mgr25__stu__ready     ),
            .stu__mgr25__type         ( stu__mgr25__type      ),
            .stu__mgr25__data         ( stu__mgr25__data      ),
            .stu__mgr25__oob_data     ( stu__mgr25__oob_data  ),

            .stu__mgr26__valid        ( stu__mgr26__valid     ),
            .stu__mgr26__cntl         ( stu__mgr26__cntl      ),
            .mgr26__stu__ready        ( mgr26__stu__ready     ),
            .stu__mgr26__type         ( stu__mgr26__type      ),
            .stu__mgr26__data         ( stu__mgr26__data      ),
            .stu__mgr26__oob_data     ( stu__mgr26__oob_data  ),

            .stu__mgr27__valid        ( stu__mgr27__valid     ),
            .stu__mgr27__cntl         ( stu__mgr27__cntl      ),
            .mgr27__stu__ready        ( mgr27__stu__ready     ),
            .stu__mgr27__type         ( stu__mgr27__type      ),
            .stu__mgr27__data         ( stu__mgr27__data      ),
            .stu__mgr27__oob_data     ( stu__mgr27__oob_data  ),

            .stu__mgr28__valid        ( stu__mgr28__valid     ),
            .stu__mgr28__cntl         ( stu__mgr28__cntl      ),
            .mgr28__stu__ready        ( mgr28__stu__ready     ),
            .stu__mgr28__type         ( stu__mgr28__type      ),
            .stu__mgr28__data         ( stu__mgr28__data      ),
            .stu__mgr28__oob_data     ( stu__mgr28__oob_data  ),

            .stu__mgr29__valid        ( stu__mgr29__valid     ),
            .stu__mgr29__cntl         ( stu__mgr29__cntl      ),
            .mgr29__stu__ready        ( mgr29__stu__ready     ),
            .stu__mgr29__type         ( stu__mgr29__type      ),
            .stu__mgr29__data         ( stu__mgr29__data      ),
            .stu__mgr29__oob_data     ( stu__mgr29__oob_data  ),

            .stu__mgr30__valid        ( stu__mgr30__valid     ),
            .stu__mgr30__cntl         ( stu__mgr30__cntl      ),
            .mgr30__stu__ready        ( mgr30__stu__ready     ),
            .stu__mgr30__type         ( stu__mgr30__type      ),
            .stu__mgr30__data         ( stu__mgr30__data      ),
            .stu__mgr30__oob_data     ( stu__mgr30__oob_data  ),

            .stu__mgr31__valid        ( stu__mgr31__valid     ),
            .stu__mgr31__cntl         ( stu__mgr31__cntl      ),
            .mgr31__stu__ready        ( mgr31__stu__ready     ),
            .stu__mgr31__type         ( stu__mgr31__type      ),
            .stu__mgr31__data         ( stu__mgr31__data      ),
            .stu__mgr31__oob_data     ( stu__mgr31__oob_data  ),

            .stu__mgr32__valid        ( stu__mgr32__valid     ),
            .stu__mgr32__cntl         ( stu__mgr32__cntl      ),
            .mgr32__stu__ready        ( mgr32__stu__ready     ),
            .stu__mgr32__type         ( stu__mgr32__type      ),
            .stu__mgr32__data         ( stu__mgr32__data      ),
            .stu__mgr32__oob_data     ( stu__mgr32__oob_data  ),

            .stu__mgr33__valid        ( stu__mgr33__valid     ),
            .stu__mgr33__cntl         ( stu__mgr33__cntl      ),
            .mgr33__stu__ready        ( mgr33__stu__ready     ),
            .stu__mgr33__type         ( stu__mgr33__type      ),
            .stu__mgr33__data         ( stu__mgr33__data      ),
            .stu__mgr33__oob_data     ( stu__mgr33__oob_data  ),

            .stu__mgr34__valid        ( stu__mgr34__valid     ),
            .stu__mgr34__cntl         ( stu__mgr34__cntl      ),
            .mgr34__stu__ready        ( mgr34__stu__ready     ),
            .stu__mgr34__type         ( stu__mgr34__type      ),
            .stu__mgr34__data         ( stu__mgr34__data      ),
            .stu__mgr34__oob_data     ( stu__mgr34__oob_data  ),

            .stu__mgr35__valid        ( stu__mgr35__valid     ),
            .stu__mgr35__cntl         ( stu__mgr35__cntl      ),
            .mgr35__stu__ready        ( mgr35__stu__ready     ),
            .stu__mgr35__type         ( stu__mgr35__type      ),
            .stu__mgr35__data         ( stu__mgr35__data      ),
            .stu__mgr35__oob_data     ( stu__mgr35__oob_data  ),

            .stu__mgr36__valid        ( stu__mgr36__valid     ),
            .stu__mgr36__cntl         ( stu__mgr36__cntl      ),
            .mgr36__stu__ready        ( mgr36__stu__ready     ),
            .stu__mgr36__type         ( stu__mgr36__type      ),
            .stu__mgr36__data         ( stu__mgr36__data      ),
            .stu__mgr36__oob_data     ( stu__mgr36__oob_data  ),

            .stu__mgr37__valid        ( stu__mgr37__valid     ),
            .stu__mgr37__cntl         ( stu__mgr37__cntl      ),
            .mgr37__stu__ready        ( mgr37__stu__ready     ),
            .stu__mgr37__type         ( stu__mgr37__type      ),
            .stu__mgr37__data         ( stu__mgr37__data      ),
            .stu__mgr37__oob_data     ( stu__mgr37__oob_data  ),

            .stu__mgr38__valid        ( stu__mgr38__valid     ),
            .stu__mgr38__cntl         ( stu__mgr38__cntl      ),
            .mgr38__stu__ready        ( mgr38__stu__ready     ),
            .stu__mgr38__type         ( stu__mgr38__type      ),
            .stu__mgr38__data         ( stu__mgr38__data      ),
            .stu__mgr38__oob_data     ( stu__mgr38__oob_data  ),

            .stu__mgr39__valid        ( stu__mgr39__valid     ),
            .stu__mgr39__cntl         ( stu__mgr39__cntl      ),
            .mgr39__stu__ready        ( mgr39__stu__ready     ),
            .stu__mgr39__type         ( stu__mgr39__type      ),
            .stu__mgr39__data         ( stu__mgr39__data      ),
            .stu__mgr39__oob_data     ( stu__mgr39__oob_data  ),

            .stu__mgr40__valid        ( stu__mgr40__valid     ),
            .stu__mgr40__cntl         ( stu__mgr40__cntl      ),
            .mgr40__stu__ready        ( mgr40__stu__ready     ),
            .stu__mgr40__type         ( stu__mgr40__type      ),
            .stu__mgr40__data         ( stu__mgr40__data      ),
            .stu__mgr40__oob_data     ( stu__mgr40__oob_data  ),

            .stu__mgr41__valid        ( stu__mgr41__valid     ),
            .stu__mgr41__cntl         ( stu__mgr41__cntl      ),
            .mgr41__stu__ready        ( mgr41__stu__ready     ),
            .stu__mgr41__type         ( stu__mgr41__type      ),
            .stu__mgr41__data         ( stu__mgr41__data      ),
            .stu__mgr41__oob_data     ( stu__mgr41__oob_data  ),

            .stu__mgr42__valid        ( stu__mgr42__valid     ),
            .stu__mgr42__cntl         ( stu__mgr42__cntl      ),
            .mgr42__stu__ready        ( mgr42__stu__ready     ),
            .stu__mgr42__type         ( stu__mgr42__type      ),
            .stu__mgr42__data         ( stu__mgr42__data      ),
            .stu__mgr42__oob_data     ( stu__mgr42__oob_data  ),

            .stu__mgr43__valid        ( stu__mgr43__valid     ),
            .stu__mgr43__cntl         ( stu__mgr43__cntl      ),
            .mgr43__stu__ready        ( mgr43__stu__ready     ),
            .stu__mgr43__type         ( stu__mgr43__type      ),
            .stu__mgr43__data         ( stu__mgr43__data      ),
            .stu__mgr43__oob_data     ( stu__mgr43__oob_data  ),

            .stu__mgr44__valid        ( stu__mgr44__valid     ),
            .stu__mgr44__cntl         ( stu__mgr44__cntl      ),
            .mgr44__stu__ready        ( mgr44__stu__ready     ),
            .stu__mgr44__type         ( stu__mgr44__type      ),
            .stu__mgr44__data         ( stu__mgr44__data      ),
            .stu__mgr44__oob_data     ( stu__mgr44__oob_data  ),

            .stu__mgr45__valid        ( stu__mgr45__valid     ),
            .stu__mgr45__cntl         ( stu__mgr45__cntl      ),
            .mgr45__stu__ready        ( mgr45__stu__ready     ),
            .stu__mgr45__type         ( stu__mgr45__type      ),
            .stu__mgr45__data         ( stu__mgr45__data      ),
            .stu__mgr45__oob_data     ( stu__mgr45__oob_data  ),

            .stu__mgr46__valid        ( stu__mgr46__valid     ),
            .stu__mgr46__cntl         ( stu__mgr46__cntl      ),
            .mgr46__stu__ready        ( mgr46__stu__ready     ),
            .stu__mgr46__type         ( stu__mgr46__type      ),
            .stu__mgr46__data         ( stu__mgr46__data      ),
            .stu__mgr46__oob_data     ( stu__mgr46__oob_data  ),

            .stu__mgr47__valid        ( stu__mgr47__valid     ),
            .stu__mgr47__cntl         ( stu__mgr47__cntl      ),
            .mgr47__stu__ready        ( mgr47__stu__ready     ),
            .stu__mgr47__type         ( stu__mgr47__type      ),
            .stu__mgr47__data         ( stu__mgr47__data      ),
            .stu__mgr47__oob_data     ( stu__mgr47__oob_data  ),

            .stu__mgr48__valid        ( stu__mgr48__valid     ),
            .stu__mgr48__cntl         ( stu__mgr48__cntl      ),
            .mgr48__stu__ready        ( mgr48__stu__ready     ),
            .stu__mgr48__type         ( stu__mgr48__type      ),
            .stu__mgr48__data         ( stu__mgr48__data      ),
            .stu__mgr48__oob_data     ( stu__mgr48__oob_data  ),

            .stu__mgr49__valid        ( stu__mgr49__valid     ),
            .stu__mgr49__cntl         ( stu__mgr49__cntl      ),
            .mgr49__stu__ready        ( mgr49__stu__ready     ),
            .stu__mgr49__type         ( stu__mgr49__type      ),
            .stu__mgr49__data         ( stu__mgr49__data      ),
            .stu__mgr49__oob_data     ( stu__mgr49__oob_data  ),

            .stu__mgr50__valid        ( stu__mgr50__valid     ),
            .stu__mgr50__cntl         ( stu__mgr50__cntl      ),
            .mgr50__stu__ready        ( mgr50__stu__ready     ),
            .stu__mgr50__type         ( stu__mgr50__type      ),
            .stu__mgr50__data         ( stu__mgr50__data      ),
            .stu__mgr50__oob_data     ( stu__mgr50__oob_data  ),

            .stu__mgr51__valid        ( stu__mgr51__valid     ),
            .stu__mgr51__cntl         ( stu__mgr51__cntl      ),
            .mgr51__stu__ready        ( mgr51__stu__ready     ),
            .stu__mgr51__type         ( stu__mgr51__type      ),
            .stu__mgr51__data         ( stu__mgr51__data      ),
            .stu__mgr51__oob_data     ( stu__mgr51__oob_data  ),

            .stu__mgr52__valid        ( stu__mgr52__valid     ),
            .stu__mgr52__cntl         ( stu__mgr52__cntl      ),
            .mgr52__stu__ready        ( mgr52__stu__ready     ),
            .stu__mgr52__type         ( stu__mgr52__type      ),
            .stu__mgr52__data         ( stu__mgr52__data      ),
            .stu__mgr52__oob_data     ( stu__mgr52__oob_data  ),

            .stu__mgr53__valid        ( stu__mgr53__valid     ),
            .stu__mgr53__cntl         ( stu__mgr53__cntl      ),
            .mgr53__stu__ready        ( mgr53__stu__ready     ),
            .stu__mgr53__type         ( stu__mgr53__type      ),
            .stu__mgr53__data         ( stu__mgr53__data      ),
            .stu__mgr53__oob_data     ( stu__mgr53__oob_data  ),

            .stu__mgr54__valid        ( stu__mgr54__valid     ),
            .stu__mgr54__cntl         ( stu__mgr54__cntl      ),
            .mgr54__stu__ready        ( mgr54__stu__ready     ),
            .stu__mgr54__type         ( stu__mgr54__type      ),
            .stu__mgr54__data         ( stu__mgr54__data      ),
            .stu__mgr54__oob_data     ( stu__mgr54__oob_data  ),

            .stu__mgr55__valid        ( stu__mgr55__valid     ),
            .stu__mgr55__cntl         ( stu__mgr55__cntl      ),
            .mgr55__stu__ready        ( mgr55__stu__ready     ),
            .stu__mgr55__type         ( stu__mgr55__type      ),
            .stu__mgr55__data         ( stu__mgr55__data      ),
            .stu__mgr55__oob_data     ( stu__mgr55__oob_data  ),

            .stu__mgr56__valid        ( stu__mgr56__valid     ),
            .stu__mgr56__cntl         ( stu__mgr56__cntl      ),
            .mgr56__stu__ready        ( mgr56__stu__ready     ),
            .stu__mgr56__type         ( stu__mgr56__type      ),
            .stu__mgr56__data         ( stu__mgr56__data      ),
            .stu__mgr56__oob_data     ( stu__mgr56__oob_data  ),

            .stu__mgr57__valid        ( stu__mgr57__valid     ),
            .stu__mgr57__cntl         ( stu__mgr57__cntl      ),
            .mgr57__stu__ready        ( mgr57__stu__ready     ),
            .stu__mgr57__type         ( stu__mgr57__type      ),
            .stu__mgr57__data         ( stu__mgr57__data      ),
            .stu__mgr57__oob_data     ( stu__mgr57__oob_data  ),

            .stu__mgr58__valid        ( stu__mgr58__valid     ),
            .stu__mgr58__cntl         ( stu__mgr58__cntl      ),
            .mgr58__stu__ready        ( mgr58__stu__ready     ),
            .stu__mgr58__type         ( stu__mgr58__type      ),
            .stu__mgr58__data         ( stu__mgr58__data      ),
            .stu__mgr58__oob_data     ( stu__mgr58__oob_data  ),

            .stu__mgr59__valid        ( stu__mgr59__valid     ),
            .stu__mgr59__cntl         ( stu__mgr59__cntl      ),
            .mgr59__stu__ready        ( mgr59__stu__ready     ),
            .stu__mgr59__type         ( stu__mgr59__type      ),
            .stu__mgr59__data         ( stu__mgr59__data      ),
            .stu__mgr59__oob_data     ( stu__mgr59__oob_data  ),

            .stu__mgr60__valid        ( stu__mgr60__valid     ),
            .stu__mgr60__cntl         ( stu__mgr60__cntl      ),
            .mgr60__stu__ready        ( mgr60__stu__ready     ),
            .stu__mgr60__type         ( stu__mgr60__type      ),
            .stu__mgr60__data         ( stu__mgr60__data      ),
            .stu__mgr60__oob_data     ( stu__mgr60__oob_data  ),

            .stu__mgr61__valid        ( stu__mgr61__valid     ),
            .stu__mgr61__cntl         ( stu__mgr61__cntl      ),
            .mgr61__stu__ready        ( mgr61__stu__ready     ),
            .stu__mgr61__type         ( stu__mgr61__type      ),
            .stu__mgr61__data         ( stu__mgr61__data      ),
            .stu__mgr61__oob_data     ( stu__mgr61__oob_data  ),

            .stu__mgr62__valid        ( stu__mgr62__valid     ),
            .stu__mgr62__cntl         ( stu__mgr62__cntl      ),
            .mgr62__stu__ready        ( mgr62__stu__ready     ),
            .stu__mgr62__type         ( stu__mgr62__type      ),
            .stu__mgr62__data         ( stu__mgr62__data      ),
            .stu__mgr62__oob_data     ( stu__mgr62__oob_data  ),

            .stu__mgr63__valid        ( stu__mgr63__valid     ),
            .stu__mgr63__cntl         ( stu__mgr63__cntl      ),
            .mgr63__stu__ready        ( mgr63__stu__ready     ),
            .stu__mgr63__type         ( stu__mgr63__type      ),
            .stu__mgr63__data         ( stu__mgr63__data      ),
            .stu__mgr63__oob_data     ( stu__mgr63__oob_data  ),

