
            // General control and status                    
            mgr0__sys__allSynchronized                    ,
            sys__mgr0__thisSynchronized                   ,
            sys__mgr0__ready                              ,
            sys__mgr0__complete                           ,

            // General control and status                    
            mgr1__sys__allSynchronized                    ,
            sys__mgr1__thisSynchronized                   ,
            sys__mgr1__ready                              ,
            sys__mgr1__complete                           ,

            // General control and status                    
            mgr2__sys__allSynchronized                    ,
            sys__mgr2__thisSynchronized                   ,
            sys__mgr2__ready                              ,
            sys__mgr2__complete                           ,

            // General control and status                    
            mgr3__sys__allSynchronized                    ,
            sys__mgr3__thisSynchronized                   ,
            sys__mgr3__ready                              ,
            sys__mgr3__complete                           ,
