
  assign  mgr0__std__oob_cntl                       =  mgr_inst[0].mgr__std__oob_cntl       ;
  assign  mgr0__std__oob_valid                      =  mgr_inst[0].mgr__std__oob_valid      ;
  assign  mgr_inst[0].std__mgr__oob_ready           =  std__mgr0__oob_ready                 ;
  assign  mgr0__std__oob_type                       =  mgr_inst[0].mgr__std__oob_type       ;
  assign  mgr0__std__oob_data                       =  mgr_inst[0].mgr__std__oob_data       ;

  assign  mgr1__std__oob_cntl                       =  mgr_inst[1].mgr__std__oob_cntl       ;
  assign  mgr1__std__oob_valid                      =  mgr_inst[1].mgr__std__oob_valid      ;
  assign  mgr_inst[1].std__mgr__oob_ready           =  std__mgr1__oob_ready                 ;
  assign  mgr1__std__oob_type                       =  mgr_inst[1].mgr__std__oob_type       ;
  assign  mgr1__std__oob_data                       =  mgr_inst[1].mgr__std__oob_data       ;

  assign  mgr2__std__oob_cntl                       =  mgr_inst[2].mgr__std__oob_cntl       ;
  assign  mgr2__std__oob_valid                      =  mgr_inst[2].mgr__std__oob_valid      ;
  assign  mgr_inst[2].std__mgr__oob_ready           =  std__mgr2__oob_ready                 ;
  assign  mgr2__std__oob_type                       =  mgr_inst[2].mgr__std__oob_type       ;
  assign  mgr2__std__oob_data                       =  mgr_inst[2].mgr__std__oob_data       ;

  assign  mgr3__std__oob_cntl                       =  mgr_inst[3].mgr__std__oob_cntl       ;
  assign  mgr3__std__oob_valid                      =  mgr_inst[3].mgr__std__oob_valid      ;
  assign  mgr_inst[3].std__mgr__oob_ready           =  std__mgr3__oob_ready                 ;
  assign  mgr3__std__oob_type                       =  mgr_inst[3].mgr__std__oob_type       ;
  assign  mgr3__std__oob_data                       =  mgr_inst[3].mgr__std__oob_data       ;

  assign  mgr4__std__oob_cntl                       =  mgr_inst[4].mgr__std__oob_cntl       ;
  assign  mgr4__std__oob_valid                      =  mgr_inst[4].mgr__std__oob_valid      ;
  assign  mgr_inst[4].std__mgr__oob_ready           =  std__mgr4__oob_ready                 ;
  assign  mgr4__std__oob_type                       =  mgr_inst[4].mgr__std__oob_type       ;
  assign  mgr4__std__oob_data                       =  mgr_inst[4].mgr__std__oob_data       ;

  assign  mgr5__std__oob_cntl                       =  mgr_inst[5].mgr__std__oob_cntl       ;
  assign  mgr5__std__oob_valid                      =  mgr_inst[5].mgr__std__oob_valid      ;
  assign  mgr_inst[5].std__mgr__oob_ready           =  std__mgr5__oob_ready                 ;
  assign  mgr5__std__oob_type                       =  mgr_inst[5].mgr__std__oob_type       ;
  assign  mgr5__std__oob_data                       =  mgr_inst[5].mgr__std__oob_data       ;

  assign  mgr6__std__oob_cntl                       =  mgr_inst[6].mgr__std__oob_cntl       ;
  assign  mgr6__std__oob_valid                      =  mgr_inst[6].mgr__std__oob_valid      ;
  assign  mgr_inst[6].std__mgr__oob_ready           =  std__mgr6__oob_ready                 ;
  assign  mgr6__std__oob_type                       =  mgr_inst[6].mgr__std__oob_type       ;
  assign  mgr6__std__oob_data                       =  mgr_inst[6].mgr__std__oob_data       ;

  assign  mgr7__std__oob_cntl                       =  mgr_inst[7].mgr__std__oob_cntl       ;
  assign  mgr7__std__oob_valid                      =  mgr_inst[7].mgr__std__oob_valid      ;
  assign  mgr_inst[7].std__mgr__oob_ready           =  std__mgr7__oob_ready                 ;
  assign  mgr7__std__oob_type                       =  mgr_inst[7].mgr__std__oob_type       ;
  assign  mgr7__std__oob_data                       =  mgr_inst[7].mgr__std__oob_data       ;

  assign  mgr8__std__oob_cntl                       =  mgr_inst[8].mgr__std__oob_cntl       ;
  assign  mgr8__std__oob_valid                      =  mgr_inst[8].mgr__std__oob_valid      ;
  assign  mgr_inst[8].std__mgr__oob_ready           =  std__mgr8__oob_ready                 ;
  assign  mgr8__std__oob_type                       =  mgr_inst[8].mgr__std__oob_type       ;
  assign  mgr8__std__oob_data                       =  mgr_inst[8].mgr__std__oob_data       ;

  assign  mgr9__std__oob_cntl                       =  mgr_inst[9].mgr__std__oob_cntl       ;
  assign  mgr9__std__oob_valid                      =  mgr_inst[9].mgr__std__oob_valid      ;
  assign  mgr_inst[9].std__mgr__oob_ready           =  std__mgr9__oob_ready                 ;
  assign  mgr9__std__oob_type                       =  mgr_inst[9].mgr__std__oob_type       ;
  assign  mgr9__std__oob_data                       =  mgr_inst[9].mgr__std__oob_data       ;

  assign  mgr10__std__oob_cntl                       =  mgr_inst[10].mgr__std__oob_cntl       ;
  assign  mgr10__std__oob_valid                      =  mgr_inst[10].mgr__std__oob_valid      ;
  assign  mgr_inst[10].std__mgr__oob_ready           =  std__mgr10__oob_ready                 ;
  assign  mgr10__std__oob_type                       =  mgr_inst[10].mgr__std__oob_type       ;
  assign  mgr10__std__oob_data                       =  mgr_inst[10].mgr__std__oob_data       ;

  assign  mgr11__std__oob_cntl                       =  mgr_inst[11].mgr__std__oob_cntl       ;
  assign  mgr11__std__oob_valid                      =  mgr_inst[11].mgr__std__oob_valid      ;
  assign  mgr_inst[11].std__mgr__oob_ready           =  std__mgr11__oob_ready                 ;
  assign  mgr11__std__oob_type                       =  mgr_inst[11].mgr__std__oob_type       ;
  assign  mgr11__std__oob_data                       =  mgr_inst[11].mgr__std__oob_data       ;

  assign  mgr12__std__oob_cntl                       =  mgr_inst[12].mgr__std__oob_cntl       ;
  assign  mgr12__std__oob_valid                      =  mgr_inst[12].mgr__std__oob_valid      ;
  assign  mgr_inst[12].std__mgr__oob_ready           =  std__mgr12__oob_ready                 ;
  assign  mgr12__std__oob_type                       =  mgr_inst[12].mgr__std__oob_type       ;
  assign  mgr12__std__oob_data                       =  mgr_inst[12].mgr__std__oob_data       ;

  assign  mgr13__std__oob_cntl                       =  mgr_inst[13].mgr__std__oob_cntl       ;
  assign  mgr13__std__oob_valid                      =  mgr_inst[13].mgr__std__oob_valid      ;
  assign  mgr_inst[13].std__mgr__oob_ready           =  std__mgr13__oob_ready                 ;
  assign  mgr13__std__oob_type                       =  mgr_inst[13].mgr__std__oob_type       ;
  assign  mgr13__std__oob_data                       =  mgr_inst[13].mgr__std__oob_data       ;

  assign  mgr14__std__oob_cntl                       =  mgr_inst[14].mgr__std__oob_cntl       ;
  assign  mgr14__std__oob_valid                      =  mgr_inst[14].mgr__std__oob_valid      ;
  assign  mgr_inst[14].std__mgr__oob_ready           =  std__mgr14__oob_ready                 ;
  assign  mgr14__std__oob_type                       =  mgr_inst[14].mgr__std__oob_type       ;
  assign  mgr14__std__oob_data                       =  mgr_inst[14].mgr__std__oob_data       ;

  assign  mgr15__std__oob_cntl                       =  mgr_inst[15].mgr__std__oob_cntl       ;
  assign  mgr15__std__oob_valid                      =  mgr_inst[15].mgr__std__oob_valid      ;
  assign  mgr_inst[15].std__mgr__oob_ready           =  std__mgr15__oob_ready                 ;
  assign  mgr15__std__oob_type                       =  mgr_inst[15].mgr__std__oob_type       ;
  assign  mgr15__std__oob_data                       =  mgr_inst[15].mgr__std__oob_data       ;

  assign  mgr16__std__oob_cntl                       =  mgr_inst[16].mgr__std__oob_cntl       ;
  assign  mgr16__std__oob_valid                      =  mgr_inst[16].mgr__std__oob_valid      ;
  assign  mgr_inst[16].std__mgr__oob_ready           =  std__mgr16__oob_ready                 ;
  assign  mgr16__std__oob_type                       =  mgr_inst[16].mgr__std__oob_type       ;
  assign  mgr16__std__oob_data                       =  mgr_inst[16].mgr__std__oob_data       ;

  assign  mgr17__std__oob_cntl                       =  mgr_inst[17].mgr__std__oob_cntl       ;
  assign  mgr17__std__oob_valid                      =  mgr_inst[17].mgr__std__oob_valid      ;
  assign  mgr_inst[17].std__mgr__oob_ready           =  std__mgr17__oob_ready                 ;
  assign  mgr17__std__oob_type                       =  mgr_inst[17].mgr__std__oob_type       ;
  assign  mgr17__std__oob_data                       =  mgr_inst[17].mgr__std__oob_data       ;

  assign  mgr18__std__oob_cntl                       =  mgr_inst[18].mgr__std__oob_cntl       ;
  assign  mgr18__std__oob_valid                      =  mgr_inst[18].mgr__std__oob_valid      ;
  assign  mgr_inst[18].std__mgr__oob_ready           =  std__mgr18__oob_ready                 ;
  assign  mgr18__std__oob_type                       =  mgr_inst[18].mgr__std__oob_type       ;
  assign  mgr18__std__oob_data                       =  mgr_inst[18].mgr__std__oob_data       ;

  assign  mgr19__std__oob_cntl                       =  mgr_inst[19].mgr__std__oob_cntl       ;
  assign  mgr19__std__oob_valid                      =  mgr_inst[19].mgr__std__oob_valid      ;
  assign  mgr_inst[19].std__mgr__oob_ready           =  std__mgr19__oob_ready                 ;
  assign  mgr19__std__oob_type                       =  mgr_inst[19].mgr__std__oob_type       ;
  assign  mgr19__std__oob_data                       =  mgr_inst[19].mgr__std__oob_data       ;

  assign  mgr20__std__oob_cntl                       =  mgr_inst[20].mgr__std__oob_cntl       ;
  assign  mgr20__std__oob_valid                      =  mgr_inst[20].mgr__std__oob_valid      ;
  assign  mgr_inst[20].std__mgr__oob_ready           =  std__mgr20__oob_ready                 ;
  assign  mgr20__std__oob_type                       =  mgr_inst[20].mgr__std__oob_type       ;
  assign  mgr20__std__oob_data                       =  mgr_inst[20].mgr__std__oob_data       ;

  assign  mgr21__std__oob_cntl                       =  mgr_inst[21].mgr__std__oob_cntl       ;
  assign  mgr21__std__oob_valid                      =  mgr_inst[21].mgr__std__oob_valid      ;
  assign  mgr_inst[21].std__mgr__oob_ready           =  std__mgr21__oob_ready                 ;
  assign  mgr21__std__oob_type                       =  mgr_inst[21].mgr__std__oob_type       ;
  assign  mgr21__std__oob_data                       =  mgr_inst[21].mgr__std__oob_data       ;

  assign  mgr22__std__oob_cntl                       =  mgr_inst[22].mgr__std__oob_cntl       ;
  assign  mgr22__std__oob_valid                      =  mgr_inst[22].mgr__std__oob_valid      ;
  assign  mgr_inst[22].std__mgr__oob_ready           =  std__mgr22__oob_ready                 ;
  assign  mgr22__std__oob_type                       =  mgr_inst[22].mgr__std__oob_type       ;
  assign  mgr22__std__oob_data                       =  mgr_inst[22].mgr__std__oob_data       ;

  assign  mgr23__std__oob_cntl                       =  mgr_inst[23].mgr__std__oob_cntl       ;
  assign  mgr23__std__oob_valid                      =  mgr_inst[23].mgr__std__oob_valid      ;
  assign  mgr_inst[23].std__mgr__oob_ready           =  std__mgr23__oob_ready                 ;
  assign  mgr23__std__oob_type                       =  mgr_inst[23].mgr__std__oob_type       ;
  assign  mgr23__std__oob_data                       =  mgr_inst[23].mgr__std__oob_data       ;

  assign  mgr24__std__oob_cntl                       =  mgr_inst[24].mgr__std__oob_cntl       ;
  assign  mgr24__std__oob_valid                      =  mgr_inst[24].mgr__std__oob_valid      ;
  assign  mgr_inst[24].std__mgr__oob_ready           =  std__mgr24__oob_ready                 ;
  assign  mgr24__std__oob_type                       =  mgr_inst[24].mgr__std__oob_type       ;
  assign  mgr24__std__oob_data                       =  mgr_inst[24].mgr__std__oob_data       ;

  assign  mgr25__std__oob_cntl                       =  mgr_inst[25].mgr__std__oob_cntl       ;
  assign  mgr25__std__oob_valid                      =  mgr_inst[25].mgr__std__oob_valid      ;
  assign  mgr_inst[25].std__mgr__oob_ready           =  std__mgr25__oob_ready                 ;
  assign  mgr25__std__oob_type                       =  mgr_inst[25].mgr__std__oob_type       ;
  assign  mgr25__std__oob_data                       =  mgr_inst[25].mgr__std__oob_data       ;

  assign  mgr26__std__oob_cntl                       =  mgr_inst[26].mgr__std__oob_cntl       ;
  assign  mgr26__std__oob_valid                      =  mgr_inst[26].mgr__std__oob_valid      ;
  assign  mgr_inst[26].std__mgr__oob_ready           =  std__mgr26__oob_ready                 ;
  assign  mgr26__std__oob_type                       =  mgr_inst[26].mgr__std__oob_type       ;
  assign  mgr26__std__oob_data                       =  mgr_inst[26].mgr__std__oob_data       ;

  assign  mgr27__std__oob_cntl                       =  mgr_inst[27].mgr__std__oob_cntl       ;
  assign  mgr27__std__oob_valid                      =  mgr_inst[27].mgr__std__oob_valid      ;
  assign  mgr_inst[27].std__mgr__oob_ready           =  std__mgr27__oob_ready                 ;
  assign  mgr27__std__oob_type                       =  mgr_inst[27].mgr__std__oob_type       ;
  assign  mgr27__std__oob_data                       =  mgr_inst[27].mgr__std__oob_data       ;

  assign  mgr28__std__oob_cntl                       =  mgr_inst[28].mgr__std__oob_cntl       ;
  assign  mgr28__std__oob_valid                      =  mgr_inst[28].mgr__std__oob_valid      ;
  assign  mgr_inst[28].std__mgr__oob_ready           =  std__mgr28__oob_ready                 ;
  assign  mgr28__std__oob_type                       =  mgr_inst[28].mgr__std__oob_type       ;
  assign  mgr28__std__oob_data                       =  mgr_inst[28].mgr__std__oob_data       ;

  assign  mgr29__std__oob_cntl                       =  mgr_inst[29].mgr__std__oob_cntl       ;
  assign  mgr29__std__oob_valid                      =  mgr_inst[29].mgr__std__oob_valid      ;
  assign  mgr_inst[29].std__mgr__oob_ready           =  std__mgr29__oob_ready                 ;
  assign  mgr29__std__oob_type                       =  mgr_inst[29].mgr__std__oob_type       ;
  assign  mgr29__std__oob_data                       =  mgr_inst[29].mgr__std__oob_data       ;

  assign  mgr30__std__oob_cntl                       =  mgr_inst[30].mgr__std__oob_cntl       ;
  assign  mgr30__std__oob_valid                      =  mgr_inst[30].mgr__std__oob_valid      ;
  assign  mgr_inst[30].std__mgr__oob_ready           =  std__mgr30__oob_ready                 ;
  assign  mgr30__std__oob_type                       =  mgr_inst[30].mgr__std__oob_type       ;
  assign  mgr30__std__oob_data                       =  mgr_inst[30].mgr__std__oob_data       ;

  assign  mgr31__std__oob_cntl                       =  mgr_inst[31].mgr__std__oob_cntl       ;
  assign  mgr31__std__oob_valid                      =  mgr_inst[31].mgr__std__oob_valid      ;
  assign  mgr_inst[31].std__mgr__oob_ready           =  std__mgr31__oob_ready                 ;
  assign  mgr31__std__oob_type                       =  mgr_inst[31].mgr__std__oob_type       ;
  assign  mgr31__std__oob_data                       =  mgr_inst[31].mgr__std__oob_data       ;

  assign  mgr32__std__oob_cntl                       =  mgr_inst[32].mgr__std__oob_cntl       ;
  assign  mgr32__std__oob_valid                      =  mgr_inst[32].mgr__std__oob_valid      ;
  assign  mgr_inst[32].std__mgr__oob_ready           =  std__mgr32__oob_ready                 ;
  assign  mgr32__std__oob_type                       =  mgr_inst[32].mgr__std__oob_type       ;
  assign  mgr32__std__oob_data                       =  mgr_inst[32].mgr__std__oob_data       ;

  assign  mgr33__std__oob_cntl                       =  mgr_inst[33].mgr__std__oob_cntl       ;
  assign  mgr33__std__oob_valid                      =  mgr_inst[33].mgr__std__oob_valid      ;
  assign  mgr_inst[33].std__mgr__oob_ready           =  std__mgr33__oob_ready                 ;
  assign  mgr33__std__oob_type                       =  mgr_inst[33].mgr__std__oob_type       ;
  assign  mgr33__std__oob_data                       =  mgr_inst[33].mgr__std__oob_data       ;

  assign  mgr34__std__oob_cntl                       =  mgr_inst[34].mgr__std__oob_cntl       ;
  assign  mgr34__std__oob_valid                      =  mgr_inst[34].mgr__std__oob_valid      ;
  assign  mgr_inst[34].std__mgr__oob_ready           =  std__mgr34__oob_ready                 ;
  assign  mgr34__std__oob_type                       =  mgr_inst[34].mgr__std__oob_type       ;
  assign  mgr34__std__oob_data                       =  mgr_inst[34].mgr__std__oob_data       ;

  assign  mgr35__std__oob_cntl                       =  mgr_inst[35].mgr__std__oob_cntl       ;
  assign  mgr35__std__oob_valid                      =  mgr_inst[35].mgr__std__oob_valid      ;
  assign  mgr_inst[35].std__mgr__oob_ready           =  std__mgr35__oob_ready                 ;
  assign  mgr35__std__oob_type                       =  mgr_inst[35].mgr__std__oob_type       ;
  assign  mgr35__std__oob_data                       =  mgr_inst[35].mgr__std__oob_data       ;

  assign  mgr36__std__oob_cntl                       =  mgr_inst[36].mgr__std__oob_cntl       ;
  assign  mgr36__std__oob_valid                      =  mgr_inst[36].mgr__std__oob_valid      ;
  assign  mgr_inst[36].std__mgr__oob_ready           =  std__mgr36__oob_ready                 ;
  assign  mgr36__std__oob_type                       =  mgr_inst[36].mgr__std__oob_type       ;
  assign  mgr36__std__oob_data                       =  mgr_inst[36].mgr__std__oob_data       ;

  assign  mgr37__std__oob_cntl                       =  mgr_inst[37].mgr__std__oob_cntl       ;
  assign  mgr37__std__oob_valid                      =  mgr_inst[37].mgr__std__oob_valid      ;
  assign  mgr_inst[37].std__mgr__oob_ready           =  std__mgr37__oob_ready                 ;
  assign  mgr37__std__oob_type                       =  mgr_inst[37].mgr__std__oob_type       ;
  assign  mgr37__std__oob_data                       =  mgr_inst[37].mgr__std__oob_data       ;

  assign  mgr38__std__oob_cntl                       =  mgr_inst[38].mgr__std__oob_cntl       ;
  assign  mgr38__std__oob_valid                      =  mgr_inst[38].mgr__std__oob_valid      ;
  assign  mgr_inst[38].std__mgr__oob_ready           =  std__mgr38__oob_ready                 ;
  assign  mgr38__std__oob_type                       =  mgr_inst[38].mgr__std__oob_type       ;
  assign  mgr38__std__oob_data                       =  mgr_inst[38].mgr__std__oob_data       ;

  assign  mgr39__std__oob_cntl                       =  mgr_inst[39].mgr__std__oob_cntl       ;
  assign  mgr39__std__oob_valid                      =  mgr_inst[39].mgr__std__oob_valid      ;
  assign  mgr_inst[39].std__mgr__oob_ready           =  std__mgr39__oob_ready                 ;
  assign  mgr39__std__oob_type                       =  mgr_inst[39].mgr__std__oob_type       ;
  assign  mgr39__std__oob_data                       =  mgr_inst[39].mgr__std__oob_data       ;

  assign  mgr40__std__oob_cntl                       =  mgr_inst[40].mgr__std__oob_cntl       ;
  assign  mgr40__std__oob_valid                      =  mgr_inst[40].mgr__std__oob_valid      ;
  assign  mgr_inst[40].std__mgr__oob_ready           =  std__mgr40__oob_ready                 ;
  assign  mgr40__std__oob_type                       =  mgr_inst[40].mgr__std__oob_type       ;
  assign  mgr40__std__oob_data                       =  mgr_inst[40].mgr__std__oob_data       ;

  assign  mgr41__std__oob_cntl                       =  mgr_inst[41].mgr__std__oob_cntl       ;
  assign  mgr41__std__oob_valid                      =  mgr_inst[41].mgr__std__oob_valid      ;
  assign  mgr_inst[41].std__mgr__oob_ready           =  std__mgr41__oob_ready                 ;
  assign  mgr41__std__oob_type                       =  mgr_inst[41].mgr__std__oob_type       ;
  assign  mgr41__std__oob_data                       =  mgr_inst[41].mgr__std__oob_data       ;

  assign  mgr42__std__oob_cntl                       =  mgr_inst[42].mgr__std__oob_cntl       ;
  assign  mgr42__std__oob_valid                      =  mgr_inst[42].mgr__std__oob_valid      ;
  assign  mgr_inst[42].std__mgr__oob_ready           =  std__mgr42__oob_ready                 ;
  assign  mgr42__std__oob_type                       =  mgr_inst[42].mgr__std__oob_type       ;
  assign  mgr42__std__oob_data                       =  mgr_inst[42].mgr__std__oob_data       ;

  assign  mgr43__std__oob_cntl                       =  mgr_inst[43].mgr__std__oob_cntl       ;
  assign  mgr43__std__oob_valid                      =  mgr_inst[43].mgr__std__oob_valid      ;
  assign  mgr_inst[43].std__mgr__oob_ready           =  std__mgr43__oob_ready                 ;
  assign  mgr43__std__oob_type                       =  mgr_inst[43].mgr__std__oob_type       ;
  assign  mgr43__std__oob_data                       =  mgr_inst[43].mgr__std__oob_data       ;

  assign  mgr44__std__oob_cntl                       =  mgr_inst[44].mgr__std__oob_cntl       ;
  assign  mgr44__std__oob_valid                      =  mgr_inst[44].mgr__std__oob_valid      ;
  assign  mgr_inst[44].std__mgr__oob_ready           =  std__mgr44__oob_ready                 ;
  assign  mgr44__std__oob_type                       =  mgr_inst[44].mgr__std__oob_type       ;
  assign  mgr44__std__oob_data                       =  mgr_inst[44].mgr__std__oob_data       ;

  assign  mgr45__std__oob_cntl                       =  mgr_inst[45].mgr__std__oob_cntl       ;
  assign  mgr45__std__oob_valid                      =  mgr_inst[45].mgr__std__oob_valid      ;
  assign  mgr_inst[45].std__mgr__oob_ready           =  std__mgr45__oob_ready                 ;
  assign  mgr45__std__oob_type                       =  mgr_inst[45].mgr__std__oob_type       ;
  assign  mgr45__std__oob_data                       =  mgr_inst[45].mgr__std__oob_data       ;

  assign  mgr46__std__oob_cntl                       =  mgr_inst[46].mgr__std__oob_cntl       ;
  assign  mgr46__std__oob_valid                      =  mgr_inst[46].mgr__std__oob_valid      ;
  assign  mgr_inst[46].std__mgr__oob_ready           =  std__mgr46__oob_ready                 ;
  assign  mgr46__std__oob_type                       =  mgr_inst[46].mgr__std__oob_type       ;
  assign  mgr46__std__oob_data                       =  mgr_inst[46].mgr__std__oob_data       ;

  assign  mgr47__std__oob_cntl                       =  mgr_inst[47].mgr__std__oob_cntl       ;
  assign  mgr47__std__oob_valid                      =  mgr_inst[47].mgr__std__oob_valid      ;
  assign  mgr_inst[47].std__mgr__oob_ready           =  std__mgr47__oob_ready                 ;
  assign  mgr47__std__oob_type                       =  mgr_inst[47].mgr__std__oob_type       ;
  assign  mgr47__std__oob_data                       =  mgr_inst[47].mgr__std__oob_data       ;

  assign  mgr48__std__oob_cntl                       =  mgr_inst[48].mgr__std__oob_cntl       ;
  assign  mgr48__std__oob_valid                      =  mgr_inst[48].mgr__std__oob_valid      ;
  assign  mgr_inst[48].std__mgr__oob_ready           =  std__mgr48__oob_ready                 ;
  assign  mgr48__std__oob_type                       =  mgr_inst[48].mgr__std__oob_type       ;
  assign  mgr48__std__oob_data                       =  mgr_inst[48].mgr__std__oob_data       ;

  assign  mgr49__std__oob_cntl                       =  mgr_inst[49].mgr__std__oob_cntl       ;
  assign  mgr49__std__oob_valid                      =  mgr_inst[49].mgr__std__oob_valid      ;
  assign  mgr_inst[49].std__mgr__oob_ready           =  std__mgr49__oob_ready                 ;
  assign  mgr49__std__oob_type                       =  mgr_inst[49].mgr__std__oob_type       ;
  assign  mgr49__std__oob_data                       =  mgr_inst[49].mgr__std__oob_data       ;

  assign  mgr50__std__oob_cntl                       =  mgr_inst[50].mgr__std__oob_cntl       ;
  assign  mgr50__std__oob_valid                      =  mgr_inst[50].mgr__std__oob_valid      ;
  assign  mgr_inst[50].std__mgr__oob_ready           =  std__mgr50__oob_ready                 ;
  assign  mgr50__std__oob_type                       =  mgr_inst[50].mgr__std__oob_type       ;
  assign  mgr50__std__oob_data                       =  mgr_inst[50].mgr__std__oob_data       ;

  assign  mgr51__std__oob_cntl                       =  mgr_inst[51].mgr__std__oob_cntl       ;
  assign  mgr51__std__oob_valid                      =  mgr_inst[51].mgr__std__oob_valid      ;
  assign  mgr_inst[51].std__mgr__oob_ready           =  std__mgr51__oob_ready                 ;
  assign  mgr51__std__oob_type                       =  mgr_inst[51].mgr__std__oob_type       ;
  assign  mgr51__std__oob_data                       =  mgr_inst[51].mgr__std__oob_data       ;

  assign  mgr52__std__oob_cntl                       =  mgr_inst[52].mgr__std__oob_cntl       ;
  assign  mgr52__std__oob_valid                      =  mgr_inst[52].mgr__std__oob_valid      ;
  assign  mgr_inst[52].std__mgr__oob_ready           =  std__mgr52__oob_ready                 ;
  assign  mgr52__std__oob_type                       =  mgr_inst[52].mgr__std__oob_type       ;
  assign  mgr52__std__oob_data                       =  mgr_inst[52].mgr__std__oob_data       ;

  assign  mgr53__std__oob_cntl                       =  mgr_inst[53].mgr__std__oob_cntl       ;
  assign  mgr53__std__oob_valid                      =  mgr_inst[53].mgr__std__oob_valid      ;
  assign  mgr_inst[53].std__mgr__oob_ready           =  std__mgr53__oob_ready                 ;
  assign  mgr53__std__oob_type                       =  mgr_inst[53].mgr__std__oob_type       ;
  assign  mgr53__std__oob_data                       =  mgr_inst[53].mgr__std__oob_data       ;

  assign  mgr54__std__oob_cntl                       =  mgr_inst[54].mgr__std__oob_cntl       ;
  assign  mgr54__std__oob_valid                      =  mgr_inst[54].mgr__std__oob_valid      ;
  assign  mgr_inst[54].std__mgr__oob_ready           =  std__mgr54__oob_ready                 ;
  assign  mgr54__std__oob_type                       =  mgr_inst[54].mgr__std__oob_type       ;
  assign  mgr54__std__oob_data                       =  mgr_inst[54].mgr__std__oob_data       ;

  assign  mgr55__std__oob_cntl                       =  mgr_inst[55].mgr__std__oob_cntl       ;
  assign  mgr55__std__oob_valid                      =  mgr_inst[55].mgr__std__oob_valid      ;
  assign  mgr_inst[55].std__mgr__oob_ready           =  std__mgr55__oob_ready                 ;
  assign  mgr55__std__oob_type                       =  mgr_inst[55].mgr__std__oob_type       ;
  assign  mgr55__std__oob_data                       =  mgr_inst[55].mgr__std__oob_data       ;

  assign  mgr56__std__oob_cntl                       =  mgr_inst[56].mgr__std__oob_cntl       ;
  assign  mgr56__std__oob_valid                      =  mgr_inst[56].mgr__std__oob_valid      ;
  assign  mgr_inst[56].std__mgr__oob_ready           =  std__mgr56__oob_ready                 ;
  assign  mgr56__std__oob_type                       =  mgr_inst[56].mgr__std__oob_type       ;
  assign  mgr56__std__oob_data                       =  mgr_inst[56].mgr__std__oob_data       ;

  assign  mgr57__std__oob_cntl                       =  mgr_inst[57].mgr__std__oob_cntl       ;
  assign  mgr57__std__oob_valid                      =  mgr_inst[57].mgr__std__oob_valid      ;
  assign  mgr_inst[57].std__mgr__oob_ready           =  std__mgr57__oob_ready                 ;
  assign  mgr57__std__oob_type                       =  mgr_inst[57].mgr__std__oob_type       ;
  assign  mgr57__std__oob_data                       =  mgr_inst[57].mgr__std__oob_data       ;

  assign  mgr58__std__oob_cntl                       =  mgr_inst[58].mgr__std__oob_cntl       ;
  assign  mgr58__std__oob_valid                      =  mgr_inst[58].mgr__std__oob_valid      ;
  assign  mgr_inst[58].std__mgr__oob_ready           =  std__mgr58__oob_ready                 ;
  assign  mgr58__std__oob_type                       =  mgr_inst[58].mgr__std__oob_type       ;
  assign  mgr58__std__oob_data                       =  mgr_inst[58].mgr__std__oob_data       ;

  assign  mgr59__std__oob_cntl                       =  mgr_inst[59].mgr__std__oob_cntl       ;
  assign  mgr59__std__oob_valid                      =  mgr_inst[59].mgr__std__oob_valid      ;
  assign  mgr_inst[59].std__mgr__oob_ready           =  std__mgr59__oob_ready                 ;
  assign  mgr59__std__oob_type                       =  mgr_inst[59].mgr__std__oob_type       ;
  assign  mgr59__std__oob_data                       =  mgr_inst[59].mgr__std__oob_data       ;

  assign  mgr60__std__oob_cntl                       =  mgr_inst[60].mgr__std__oob_cntl       ;
  assign  mgr60__std__oob_valid                      =  mgr_inst[60].mgr__std__oob_valid      ;
  assign  mgr_inst[60].std__mgr__oob_ready           =  std__mgr60__oob_ready                 ;
  assign  mgr60__std__oob_type                       =  mgr_inst[60].mgr__std__oob_type       ;
  assign  mgr60__std__oob_data                       =  mgr_inst[60].mgr__std__oob_data       ;

  assign  mgr61__std__oob_cntl                       =  mgr_inst[61].mgr__std__oob_cntl       ;
  assign  mgr61__std__oob_valid                      =  mgr_inst[61].mgr__std__oob_valid      ;
  assign  mgr_inst[61].std__mgr__oob_ready           =  std__mgr61__oob_ready                 ;
  assign  mgr61__std__oob_type                       =  mgr_inst[61].mgr__std__oob_type       ;
  assign  mgr61__std__oob_data                       =  mgr_inst[61].mgr__std__oob_data       ;

  assign  mgr62__std__oob_cntl                       =  mgr_inst[62].mgr__std__oob_cntl       ;
  assign  mgr62__std__oob_valid                      =  mgr_inst[62].mgr__std__oob_valid      ;
  assign  mgr_inst[62].std__mgr__oob_ready           =  std__mgr62__oob_ready                 ;
  assign  mgr62__std__oob_type                       =  mgr_inst[62].mgr__std__oob_type       ;
  assign  mgr62__std__oob_data                       =  mgr_inst[62].mgr__std__oob_data       ;

  assign  mgr63__std__oob_cntl                       =  mgr_inst[63].mgr__std__oob_cntl       ;
  assign  mgr63__std__oob_valid                      =  mgr_inst[63].mgr__std__oob_valid      ;
  assign  mgr_inst[63].std__mgr__oob_ready           =  std__mgr63__oob_ready                 ;
  assign  mgr63__std__oob_type                       =  mgr_inst[63].mgr__std__oob_type       ;
  assign  mgr63__std__oob_data                       =  mgr_inst[63].mgr__std__oob_data       ;

