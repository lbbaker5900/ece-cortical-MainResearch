
  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      mgr0__std__oob_cntl            ;
  wire                                        mgr0__std__oob_valid           ;
  wire                                        std__mgr0__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr0__std__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr0__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      mgr1__std__oob_cntl            ;
  wire                                        mgr1__std__oob_valid           ;
  wire                                        std__mgr1__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr1__std__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr1__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      mgr2__std__oob_cntl            ;
  wire                                        mgr2__std__oob_valid           ;
  wire                                        std__mgr2__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr2__std__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr2__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                
  wire[`COMMON_STD_INTF_CNTL_RANGE     ]      mgr3__std__oob_cntl            ;
  wire                                        mgr3__std__oob_valid           ;
  wire                                        std__mgr3__oob_ready           ;
  wire[`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr3__std__oob_type            ;
  wire[`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr3__std__oob_data            ;
