
            begin
              mr_proc[0][0].run()  ;
            end

            begin
              mr_proc[0][1].run()  ;
            end

            begin
              mr_proc[1][0].run()  ;
            end

            begin
              mr_proc[1][1].run()  ;
            end

            begin
              mr_proc[2][0].run()  ;
            end

            begin
              mr_proc[2][1].run()  ;
            end

            begin
              mr_proc[3][0].run()  ;
            end

            begin
              mr_proc[3][1].run()  ;
            end

            begin
              mr_proc[4][0].run()  ;
            end

            begin
              mr_proc[4][1].run()  ;
            end

            begin
              mr_proc[5][0].run()  ;
            end

            begin
              mr_proc[5][1].run()  ;
            end

            begin
              mr_proc[6][0].run()  ;
            end

            begin
              mr_proc[6][1].run()  ;
            end

            begin
              mr_proc[7][0].run()  ;
            end

            begin
              mr_proc[7][1].run()  ;
            end

            begin
              mr_proc[8][0].run()  ;
            end

            begin
              mr_proc[8][1].run()  ;
            end

            begin
              mr_proc[9][0].run()  ;
            end

            begin
              mr_proc[9][1].run()  ;
            end

            begin
              mr_proc[10][0].run()  ;
            end

            begin
              mr_proc[10][1].run()  ;
            end

            begin
              mr_proc[11][0].run()  ;
            end

            begin
              mr_proc[11][1].run()  ;
            end

            begin
              mr_proc[12][0].run()  ;
            end

            begin
              mr_proc[12][1].run()  ;
            end

            begin
              mr_proc[13][0].run()  ;
            end

            begin
              mr_proc[13][1].run()  ;
            end

            begin
              mr_proc[14][0].run()  ;
            end

            begin
              mr_proc[14][1].run()  ;
            end

            begin
              mr_proc[15][0].run()  ;
            end

            begin
              mr_proc[15][1].run()  ;
            end

            begin
              mr_proc[16][0].run()  ;
            end

            begin
              mr_proc[16][1].run()  ;
            end

            begin
              mr_proc[17][0].run()  ;
            end

            begin
              mr_proc[17][1].run()  ;
            end

            begin
              mr_proc[18][0].run()  ;
            end

            begin
              mr_proc[18][1].run()  ;
            end

            begin
              mr_proc[19][0].run()  ;
            end

            begin
              mr_proc[19][1].run()  ;
            end

            begin
              mr_proc[20][0].run()  ;
            end

            begin
              mr_proc[20][1].run()  ;
            end

            begin
              mr_proc[21][0].run()  ;
            end

            begin
              mr_proc[21][1].run()  ;
            end

            begin
              mr_proc[22][0].run()  ;
            end

            begin
              mr_proc[22][1].run()  ;
            end

            begin
              mr_proc[23][0].run()  ;
            end

            begin
              mr_proc[23][1].run()  ;
            end

            begin
              mr_proc[24][0].run()  ;
            end

            begin
              mr_proc[24][1].run()  ;
            end

            begin
              mr_proc[25][0].run()  ;
            end

            begin
              mr_proc[25][1].run()  ;
            end

            begin
              mr_proc[26][0].run()  ;
            end

            begin
              mr_proc[26][1].run()  ;
            end

            begin
              mr_proc[27][0].run()  ;
            end

            begin
              mr_proc[27][1].run()  ;
            end

            begin
              mr_proc[28][0].run()  ;
            end

            begin
              mr_proc[28][1].run()  ;
            end

            begin
              mr_proc[29][0].run()  ;
            end

            begin
              mr_proc[29][1].run()  ;
            end

            begin
              mr_proc[30][0].run()  ;
            end

            begin
              mr_proc[30][1].run()  ;
            end

            begin
              mr_proc[31][0].run()  ;
            end

            begin
              mr_proc[31][1].run()  ;
            end

            begin
              mr_proc[32][0].run()  ;
            end

            begin
              mr_proc[32][1].run()  ;
            end

            begin
              mr_proc[33][0].run()  ;
            end

            begin
              mr_proc[33][1].run()  ;
            end

            begin
              mr_proc[34][0].run()  ;
            end

            begin
              mr_proc[34][1].run()  ;
            end

            begin
              mr_proc[35][0].run()  ;
            end

            begin
              mr_proc[35][1].run()  ;
            end

            begin
              mr_proc[36][0].run()  ;
            end

            begin
              mr_proc[36][1].run()  ;
            end

            begin
              mr_proc[37][0].run()  ;
            end

            begin
              mr_proc[37][1].run()  ;
            end

            begin
              mr_proc[38][0].run()  ;
            end

            begin
              mr_proc[38][1].run()  ;
            end

            begin
              mr_proc[39][0].run()  ;
            end

            begin
              mr_proc[39][1].run()  ;
            end

            begin
              mr_proc[40][0].run()  ;
            end

            begin
              mr_proc[40][1].run()  ;
            end

            begin
              mr_proc[41][0].run()  ;
            end

            begin
              mr_proc[41][1].run()  ;
            end

            begin
              mr_proc[42][0].run()  ;
            end

            begin
              mr_proc[42][1].run()  ;
            end

            begin
              mr_proc[43][0].run()  ;
            end

            begin
              mr_proc[43][1].run()  ;
            end

            begin
              mr_proc[44][0].run()  ;
            end

            begin
              mr_proc[44][1].run()  ;
            end

            begin
              mr_proc[45][0].run()  ;
            end

            begin
              mr_proc[45][1].run()  ;
            end

            begin
              mr_proc[46][0].run()  ;
            end

            begin
              mr_proc[46][1].run()  ;
            end

            begin
              mr_proc[47][0].run()  ;
            end

            begin
              mr_proc[47][1].run()  ;
            end

            begin
              mr_proc[48][0].run()  ;
            end

            begin
              mr_proc[48][1].run()  ;
            end

            begin
              mr_proc[49][0].run()  ;
            end

            begin
              mr_proc[49][1].run()  ;
            end

            begin
              mr_proc[50][0].run()  ;
            end

            begin
              mr_proc[50][1].run()  ;
            end

            begin
              mr_proc[51][0].run()  ;
            end

            begin
              mr_proc[51][1].run()  ;
            end

            begin
              mr_proc[52][0].run()  ;
            end

            begin
              mr_proc[52][1].run()  ;
            end

            begin
              mr_proc[53][0].run()  ;
            end

            begin
              mr_proc[53][1].run()  ;
            end

            begin
              mr_proc[54][0].run()  ;
            end

            begin
              mr_proc[54][1].run()  ;
            end

            begin
              mr_proc[55][0].run()  ;
            end

            begin
              mr_proc[55][1].run()  ;
            end

            begin
              mr_proc[56][0].run()  ;
            end

            begin
              mr_proc[56][1].run()  ;
            end

            begin
              mr_proc[57][0].run()  ;
            end

            begin
              mr_proc[57][1].run()  ;
            end

            begin
              mr_proc[58][0].run()  ;
            end

            begin
              mr_proc[58][1].run()  ;
            end

            begin
              mr_proc[59][0].run()  ;
            end

            begin
              mr_proc[59][1].run()  ;
            end

            begin
              mr_proc[60][0].run()  ;
            end

            begin
              mr_proc[60][1].run()  ;
            end

            begin
              mr_proc[61][0].run()  ;
            end

            begin
              mr_proc[61][1].run()  ;
            end

            begin
              mr_proc[62][0].run()  ;
            end

            begin
              mr_proc[62][1].run()  ;
            end

            begin
              mr_proc[63][0].run()  ;
            end

            begin
              mr_proc[63][1].run()  ;
            end
