
  wire                                    reg__scntl__lane0_ready    ;
  reg                                     scntl__reg__lane0_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane0_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane0_data     ;

  wire                                    reg__scntl__lane1_ready    ;
  reg                                     scntl__reg__lane1_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane1_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane1_data     ;

  wire                                    reg__scntl__lane2_ready    ;
  reg                                     scntl__reg__lane2_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane2_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane2_data     ;

  wire                                    reg__scntl__lane3_ready    ;
  reg                                     scntl__reg__lane3_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane3_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane3_data     ;

  wire                                    reg__scntl__lane4_ready    ;
  reg                                     scntl__reg__lane4_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane4_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane4_data     ;

  wire                                    reg__scntl__lane5_ready    ;
  reg                                     scntl__reg__lane5_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane5_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane5_data     ;

  wire                                    reg__scntl__lane6_ready    ;
  reg                                     scntl__reg__lane6_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane6_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane6_data     ;

  wire                                    reg__scntl__lane7_ready    ;
  reg                                     scntl__reg__lane7_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane7_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane7_data     ;

  wire                                    reg__scntl__lane8_ready    ;
  reg                                     scntl__reg__lane8_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane8_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane8_data     ;

  wire                                    reg__scntl__lane9_ready    ;
  reg                                     scntl__reg__lane9_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane9_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane9_data     ;

  wire                                    reg__scntl__lane10_ready    ;
  reg                                     scntl__reg__lane10_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane10_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane10_data     ;

  wire                                    reg__scntl__lane11_ready    ;
  reg                                     scntl__reg__lane11_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane11_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane11_data     ;

  wire                                    reg__scntl__lane12_ready    ;
  reg                                     scntl__reg__lane12_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane12_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane12_data     ;

  wire                                    reg__scntl__lane13_ready    ;
  reg                                     scntl__reg__lane13_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane13_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane13_data     ;

  wire                                    reg__scntl__lane14_ready    ;
  reg                                     scntl__reg__lane14_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane14_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane14_data     ;

  wire                                    reg__scntl__lane15_ready    ;
  reg                                     scntl__reg__lane15_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane15_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane15_data     ;

  wire                                    reg__scntl__lane16_ready    ;
  reg                                     scntl__reg__lane16_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane16_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane16_data     ;

  wire                                    reg__scntl__lane17_ready    ;
  reg                                     scntl__reg__lane17_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane17_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane17_data     ;

  wire                                    reg__scntl__lane18_ready    ;
  reg                                     scntl__reg__lane18_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane18_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane18_data     ;

  wire                                    reg__scntl__lane19_ready    ;
  reg                                     scntl__reg__lane19_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane19_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane19_data     ;

  wire                                    reg__scntl__lane20_ready    ;
  reg                                     scntl__reg__lane20_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane20_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane20_data     ;

  wire                                    reg__scntl__lane21_ready    ;
  reg                                     scntl__reg__lane21_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane21_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane21_data     ;

  wire                                    reg__scntl__lane22_ready    ;
  reg                                     scntl__reg__lane22_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane22_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane22_data     ;

  wire                                    reg__scntl__lane23_ready    ;
  reg                                     scntl__reg__lane23_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane23_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane23_data     ;

  wire                                    reg__scntl__lane24_ready    ;
  reg                                     scntl__reg__lane24_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane24_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane24_data     ;

  wire                                    reg__scntl__lane25_ready    ;
  reg                                     scntl__reg__lane25_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane25_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane25_data     ;

  wire                                    reg__scntl__lane26_ready    ;
  reg                                     scntl__reg__lane26_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane26_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane26_data     ;

  wire                                    reg__scntl__lane27_ready    ;
  reg                                     scntl__reg__lane27_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane27_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane27_data     ;

  wire                                    reg__scntl__lane28_ready    ;
  reg                                     scntl__reg__lane28_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane28_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane28_data     ;

  wire                                    reg__scntl__lane29_ready    ;
  reg                                     scntl__reg__lane29_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane29_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane29_data     ;

  wire                                    reg__scntl__lane30_ready    ;
  reg                                     scntl__reg__lane30_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane30_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane30_data     ;

  wire                                    reg__scntl__lane31_ready    ;
  reg                                     scntl__reg__lane31_valid    ;
  reg    [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane31_cntl     ;
  reg    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane31_data     ;

