
               // General control and status                                                 
               .sys__mgr__mgrId                     ( sys__mgr__mgrId                  ),      
               .mgr__sys__allSynchronized           ( mgr__sys__allSynchronized        ),      
               .sys__mgr__thisSynchronized          ( sys__mgr__thisSynchronized       ),      
               .sys__mgr__ready                     ( sys__mgr__ready                  ),      
               .sys__mgr__complete                  ( sys__mgr__complete               ),      