
    // Common (Scalar) Register(s)                
            simd__scntl__rs0                  ,
            simd__scntl__rs1                  ,

    // Lane Registers                 
            simd__scntl__lane_r128                  ,
            simd__scntl__lane_r129                  ,
            simd__scntl__lane_r130                  ,
            simd__scntl__lane_r131                  ,
            simd__scntl__lane_r132                  ,
            simd__scntl__lane_r133                  ,
            simd__scntl__lane_r134                  ,
            simd__scntl__lane_r135                  ,
