
    // PE0, Port0 next hop mask                 
    assign pe_inst[0].sys__pe__port0_destinationMask    = `NOC_CONT_PE0_PORT0_DESTINATION_PE_BITMASK ;
    // PE0, Port1 next hop mask                 
    assign pe_inst[0].sys__pe__port1_destinationMask    = `NOC_CONT_PE0_PORT1_DESTINATION_PE_BITMASK ;
    // PE0, Port2 next hop mask                 
    assign pe_inst[0].sys__pe__port2_destinationMask    = `NOC_CONT_PE0_PORT2_DESTINATION_PE_BITMASK ;
    // PE0, Port3 next hop mask                 
    assign pe_inst[0].sys__pe__port3_destinationMask    = `NOC_CONT_PE0_PORT3_DESTINATION_PE_BITMASK ;
    // PE1, Port0 next hop mask                 
    assign pe_inst[1].sys__pe__port0_destinationMask    = `NOC_CONT_PE1_PORT0_DESTINATION_PE_BITMASK ;
    // PE1, Port1 next hop mask                 
    assign pe_inst[1].sys__pe__port1_destinationMask    = `NOC_CONT_PE1_PORT1_DESTINATION_PE_BITMASK ;
    // PE1, Port2 next hop mask                 
    assign pe_inst[1].sys__pe__port2_destinationMask    = `NOC_CONT_PE1_PORT2_DESTINATION_PE_BITMASK ;
    // PE1, Port3 next hop mask                 
    assign pe_inst[1].sys__pe__port3_destinationMask    = `NOC_CONT_PE1_PORT3_DESTINATION_PE_BITMASK ;
    // PE2, Port0 next hop mask                 
    assign pe_inst[2].sys__pe__port0_destinationMask    = `NOC_CONT_PE2_PORT0_DESTINATION_PE_BITMASK ;
    // PE2, Port1 next hop mask                 
    assign pe_inst[2].sys__pe__port1_destinationMask    = `NOC_CONT_PE2_PORT1_DESTINATION_PE_BITMASK ;
    // PE2, Port2 next hop mask                 
    assign pe_inst[2].sys__pe__port2_destinationMask    = `NOC_CONT_PE2_PORT2_DESTINATION_PE_BITMASK ;
    // PE2, Port3 next hop mask                 
    assign pe_inst[2].sys__pe__port3_destinationMask    = `NOC_CONT_PE2_PORT3_DESTINATION_PE_BITMASK ;
    // PE3, Port0 next hop mask                 
    assign pe_inst[3].sys__pe__port0_destinationMask    = `NOC_CONT_PE3_PORT0_DESTINATION_PE_BITMASK ;
    // PE3, Port1 next hop mask                 
    assign pe_inst[3].sys__pe__port1_destinationMask    = `NOC_CONT_PE3_PORT1_DESTINATION_PE_BITMASK ;
    // PE3, Port2 next hop mask                 
    assign pe_inst[3].sys__pe__port2_destinationMask    = `NOC_CONT_PE3_PORT2_DESTINATION_PE_BITMASK ;
    // PE3, Port3 next hop mask                 
    assign pe_inst[3].sys__pe__port3_destinationMask    = `NOC_CONT_PE3_PORT3_DESTINATION_PE_BITMASK ;