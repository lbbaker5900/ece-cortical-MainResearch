
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[0].put(sys_operation_lane_gen[0])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[0];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[1].put(sys_operation_lane_gen[1])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[1];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[2].put(sys_operation_lane_gen[2])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[2];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[3].put(sys_operation_lane_gen[3])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[3];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[4].put(sys_operation_lane_gen[4])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[4];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[5].put(sys_operation_lane_gen[5])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[5];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[6].put(sys_operation_lane_gen[6])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[6];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[7].put(sys_operation_lane_gen[7])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[7];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[8].put(sys_operation_lane_gen[8])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[8];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[9].put(sys_operation_lane_gen[9])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[9];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[10].put(sys_operation_lane_gen[10])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[10];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[11].put(sys_operation_lane_gen[11])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[11];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[12].put(sys_operation_lane_gen[12])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[12];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[13].put(sys_operation_lane_gen[13])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[13];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[14].put(sys_operation_lane_gen[14])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[14];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[15].put(sys_operation_lane_gen[15])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[15];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[16].put(sys_operation_lane_gen[16])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[16];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[17].put(sys_operation_lane_gen[17])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[17];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[18].put(sys_operation_lane_gen[18])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[18];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[19].put(sys_operation_lane_gen[19])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[19];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[20].put(sys_operation_lane_gen[20])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[20];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[21].put(sys_operation_lane_gen[21])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[21];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[22].put(sys_operation_lane_gen[22])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[22];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[23].put(sys_operation_lane_gen[23])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[23];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[24].put(sys_operation_lane_gen[24])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[24];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[25].put(sys_operation_lane_gen[25])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[25];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[26].put(sys_operation_lane_gen[26])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[26];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[27].put(sys_operation_lane_gen[27])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[27];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[28].put(sys_operation_lane_gen[28])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[28];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[29].put(sys_operation_lane_gen[29])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[29];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[30].put(sys_operation_lane_gen[30])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[30];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
            fork                                                                                                                                  

                // Send to driver                                                                                                                 
                mgr2gen[31].put(sys_operation_lane_gen[31])                    ;                                                                
                                                                                                                                                  
                // now wait for generator                                                                                                         
                @mgr2gen_ack[31];                                                                                                                
                                                                                                                                                  
            join_none                                                                                                                             
                                                                                                                                                  
