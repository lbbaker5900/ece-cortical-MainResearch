
  assign stOp_lane[0].cntl__stOp__operation    = cntl__sdp__lane0_stOp_operation   ;
  assign stOp_lane[0].cntl__stOp__strm0_source       = cntl__sdp__lane0_strm0_stOp_source      ;
  assign stOp_lane[0].cntl__stOp__strm0_destination  = cntl__sdp__lane0_strm0_stOp_destination ;
  assign stOp_lane[0].cntl__stOp__strm1_source       = cntl__sdp__lane0_strm1_stOp_source      ;
  assign stOp_lane[0].cntl__stOp__strm1_destination  = cntl__sdp__lane0_strm1_stOp_destination ;
  assign stOp_lane[0].cntl__stOp__strm0_enable       = cntl__sdp__lane0_strm0_stOp_enable      ;
  assign sdp__cntl__lane0_strm0_stOp_ready           = stOp_lane[0].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane0_strm0_stOp_complete        = stOp_lane[0].stOp__cntl__strm0_complete ;
  assign stOp_lane[0].cntl__stOp__strm1_enable       = cntl__sdp__lane0_strm1_stOp_enable      ;
  assign sdp__cntl__lane0_strm1_stOp_ready           = stOp_lane[0].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane0_strm1_stOp_complete        = stOp_lane[0].stOp__cntl__strm1_complete ;
  assign stOp_lane[1].cntl__stOp__operation    = cntl__sdp__lane1_stOp_operation   ;
  assign stOp_lane[1].cntl__stOp__strm0_source       = cntl__sdp__lane1_strm0_stOp_source      ;
  assign stOp_lane[1].cntl__stOp__strm0_destination  = cntl__sdp__lane1_strm0_stOp_destination ;
  assign stOp_lane[1].cntl__stOp__strm1_source       = cntl__sdp__lane1_strm1_stOp_source      ;
  assign stOp_lane[1].cntl__stOp__strm1_destination  = cntl__sdp__lane1_strm1_stOp_destination ;
  assign stOp_lane[1].cntl__stOp__strm0_enable       = cntl__sdp__lane1_strm0_stOp_enable      ;
  assign sdp__cntl__lane1_strm0_stOp_ready           = stOp_lane[1].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane1_strm0_stOp_complete        = stOp_lane[1].stOp__cntl__strm0_complete ;
  assign stOp_lane[1].cntl__stOp__strm1_enable       = cntl__sdp__lane1_strm1_stOp_enable      ;
  assign sdp__cntl__lane1_strm1_stOp_ready           = stOp_lane[1].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane1_strm1_stOp_complete        = stOp_lane[1].stOp__cntl__strm1_complete ;
  assign stOp_lane[2].cntl__stOp__operation    = cntl__sdp__lane2_stOp_operation   ;
  assign stOp_lane[2].cntl__stOp__strm0_source       = cntl__sdp__lane2_strm0_stOp_source      ;
  assign stOp_lane[2].cntl__stOp__strm0_destination  = cntl__sdp__lane2_strm0_stOp_destination ;
  assign stOp_lane[2].cntl__stOp__strm1_source       = cntl__sdp__lane2_strm1_stOp_source      ;
  assign stOp_lane[2].cntl__stOp__strm1_destination  = cntl__sdp__lane2_strm1_stOp_destination ;
  assign stOp_lane[2].cntl__stOp__strm0_enable       = cntl__sdp__lane2_strm0_stOp_enable      ;
  assign sdp__cntl__lane2_strm0_stOp_ready           = stOp_lane[2].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane2_strm0_stOp_complete        = stOp_lane[2].stOp__cntl__strm0_complete ;
  assign stOp_lane[2].cntl__stOp__strm1_enable       = cntl__sdp__lane2_strm1_stOp_enable      ;
  assign sdp__cntl__lane2_strm1_stOp_ready           = stOp_lane[2].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane2_strm1_stOp_complete        = stOp_lane[2].stOp__cntl__strm1_complete ;
  assign stOp_lane[3].cntl__stOp__operation    = cntl__sdp__lane3_stOp_operation   ;
  assign stOp_lane[3].cntl__stOp__strm0_source       = cntl__sdp__lane3_strm0_stOp_source      ;
  assign stOp_lane[3].cntl__stOp__strm0_destination  = cntl__sdp__lane3_strm0_stOp_destination ;
  assign stOp_lane[3].cntl__stOp__strm1_source       = cntl__sdp__lane3_strm1_stOp_source      ;
  assign stOp_lane[3].cntl__stOp__strm1_destination  = cntl__sdp__lane3_strm1_stOp_destination ;
  assign stOp_lane[3].cntl__stOp__strm0_enable       = cntl__sdp__lane3_strm0_stOp_enable      ;
  assign sdp__cntl__lane3_strm0_stOp_ready           = stOp_lane[3].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane3_strm0_stOp_complete        = stOp_lane[3].stOp__cntl__strm0_complete ;
  assign stOp_lane[3].cntl__stOp__strm1_enable       = cntl__sdp__lane3_strm1_stOp_enable      ;
  assign sdp__cntl__lane3_strm1_stOp_ready           = stOp_lane[3].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane3_strm1_stOp_complete        = stOp_lane[3].stOp__cntl__strm1_complete ;
  assign stOp_lane[4].cntl__stOp__operation    = cntl__sdp__lane4_stOp_operation   ;
  assign stOp_lane[4].cntl__stOp__strm0_source       = cntl__sdp__lane4_strm0_stOp_source      ;
  assign stOp_lane[4].cntl__stOp__strm0_destination  = cntl__sdp__lane4_strm0_stOp_destination ;
  assign stOp_lane[4].cntl__stOp__strm1_source       = cntl__sdp__lane4_strm1_stOp_source      ;
  assign stOp_lane[4].cntl__stOp__strm1_destination  = cntl__sdp__lane4_strm1_stOp_destination ;
  assign stOp_lane[4].cntl__stOp__strm0_enable       = cntl__sdp__lane4_strm0_stOp_enable      ;
  assign sdp__cntl__lane4_strm0_stOp_ready           = stOp_lane[4].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane4_strm0_stOp_complete        = stOp_lane[4].stOp__cntl__strm0_complete ;
  assign stOp_lane[4].cntl__stOp__strm1_enable       = cntl__sdp__lane4_strm1_stOp_enable      ;
  assign sdp__cntl__lane4_strm1_stOp_ready           = stOp_lane[4].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane4_strm1_stOp_complete        = stOp_lane[4].stOp__cntl__strm1_complete ;
  assign stOp_lane[5].cntl__stOp__operation    = cntl__sdp__lane5_stOp_operation   ;
  assign stOp_lane[5].cntl__stOp__strm0_source       = cntl__sdp__lane5_strm0_stOp_source      ;
  assign stOp_lane[5].cntl__stOp__strm0_destination  = cntl__sdp__lane5_strm0_stOp_destination ;
  assign stOp_lane[5].cntl__stOp__strm1_source       = cntl__sdp__lane5_strm1_stOp_source      ;
  assign stOp_lane[5].cntl__stOp__strm1_destination  = cntl__sdp__lane5_strm1_stOp_destination ;
  assign stOp_lane[5].cntl__stOp__strm0_enable       = cntl__sdp__lane5_strm0_stOp_enable      ;
  assign sdp__cntl__lane5_strm0_stOp_ready           = stOp_lane[5].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane5_strm0_stOp_complete        = stOp_lane[5].stOp__cntl__strm0_complete ;
  assign stOp_lane[5].cntl__stOp__strm1_enable       = cntl__sdp__lane5_strm1_stOp_enable      ;
  assign sdp__cntl__lane5_strm1_stOp_ready           = stOp_lane[5].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane5_strm1_stOp_complete        = stOp_lane[5].stOp__cntl__strm1_complete ;
  assign stOp_lane[6].cntl__stOp__operation    = cntl__sdp__lane6_stOp_operation   ;
  assign stOp_lane[6].cntl__stOp__strm0_source       = cntl__sdp__lane6_strm0_stOp_source      ;
  assign stOp_lane[6].cntl__stOp__strm0_destination  = cntl__sdp__lane6_strm0_stOp_destination ;
  assign stOp_lane[6].cntl__stOp__strm1_source       = cntl__sdp__lane6_strm1_stOp_source      ;
  assign stOp_lane[6].cntl__stOp__strm1_destination  = cntl__sdp__lane6_strm1_stOp_destination ;
  assign stOp_lane[6].cntl__stOp__strm0_enable       = cntl__sdp__lane6_strm0_stOp_enable      ;
  assign sdp__cntl__lane6_strm0_stOp_ready           = stOp_lane[6].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane6_strm0_stOp_complete        = stOp_lane[6].stOp__cntl__strm0_complete ;
  assign stOp_lane[6].cntl__stOp__strm1_enable       = cntl__sdp__lane6_strm1_stOp_enable      ;
  assign sdp__cntl__lane6_strm1_stOp_ready           = stOp_lane[6].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane6_strm1_stOp_complete        = stOp_lane[6].stOp__cntl__strm1_complete ;
  assign stOp_lane[7].cntl__stOp__operation    = cntl__sdp__lane7_stOp_operation   ;
  assign stOp_lane[7].cntl__stOp__strm0_source       = cntl__sdp__lane7_strm0_stOp_source      ;
  assign stOp_lane[7].cntl__stOp__strm0_destination  = cntl__sdp__lane7_strm0_stOp_destination ;
  assign stOp_lane[7].cntl__stOp__strm1_source       = cntl__sdp__lane7_strm1_stOp_source      ;
  assign stOp_lane[7].cntl__stOp__strm1_destination  = cntl__sdp__lane7_strm1_stOp_destination ;
  assign stOp_lane[7].cntl__stOp__strm0_enable       = cntl__sdp__lane7_strm0_stOp_enable      ;
  assign sdp__cntl__lane7_strm0_stOp_ready           = stOp_lane[7].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane7_strm0_stOp_complete        = stOp_lane[7].stOp__cntl__strm0_complete ;
  assign stOp_lane[7].cntl__stOp__strm1_enable       = cntl__sdp__lane7_strm1_stOp_enable      ;
  assign sdp__cntl__lane7_strm1_stOp_ready           = stOp_lane[7].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane7_strm1_stOp_complete        = stOp_lane[7].stOp__cntl__strm1_complete ;
  assign stOp_lane[8].cntl__stOp__operation    = cntl__sdp__lane8_stOp_operation   ;
  assign stOp_lane[8].cntl__stOp__strm0_source       = cntl__sdp__lane8_strm0_stOp_source      ;
  assign stOp_lane[8].cntl__stOp__strm0_destination  = cntl__sdp__lane8_strm0_stOp_destination ;
  assign stOp_lane[8].cntl__stOp__strm1_source       = cntl__sdp__lane8_strm1_stOp_source      ;
  assign stOp_lane[8].cntl__stOp__strm1_destination  = cntl__sdp__lane8_strm1_stOp_destination ;
  assign stOp_lane[8].cntl__stOp__strm0_enable       = cntl__sdp__lane8_strm0_stOp_enable      ;
  assign sdp__cntl__lane8_strm0_stOp_ready           = stOp_lane[8].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane8_strm0_stOp_complete        = stOp_lane[8].stOp__cntl__strm0_complete ;
  assign stOp_lane[8].cntl__stOp__strm1_enable       = cntl__sdp__lane8_strm1_stOp_enable      ;
  assign sdp__cntl__lane8_strm1_stOp_ready           = stOp_lane[8].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane8_strm1_stOp_complete        = stOp_lane[8].stOp__cntl__strm1_complete ;
  assign stOp_lane[9].cntl__stOp__operation    = cntl__sdp__lane9_stOp_operation   ;
  assign stOp_lane[9].cntl__stOp__strm0_source       = cntl__sdp__lane9_strm0_stOp_source      ;
  assign stOp_lane[9].cntl__stOp__strm0_destination  = cntl__sdp__lane9_strm0_stOp_destination ;
  assign stOp_lane[9].cntl__stOp__strm1_source       = cntl__sdp__lane9_strm1_stOp_source      ;
  assign stOp_lane[9].cntl__stOp__strm1_destination  = cntl__sdp__lane9_strm1_stOp_destination ;
  assign stOp_lane[9].cntl__stOp__strm0_enable       = cntl__sdp__lane9_strm0_stOp_enable      ;
  assign sdp__cntl__lane9_strm0_stOp_ready           = stOp_lane[9].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane9_strm0_stOp_complete        = stOp_lane[9].stOp__cntl__strm0_complete ;
  assign stOp_lane[9].cntl__stOp__strm1_enable       = cntl__sdp__lane9_strm1_stOp_enable      ;
  assign sdp__cntl__lane9_strm1_stOp_ready           = stOp_lane[9].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane9_strm1_stOp_complete        = stOp_lane[9].stOp__cntl__strm1_complete ;
  assign stOp_lane[10].cntl__stOp__operation    = cntl__sdp__lane10_stOp_operation   ;
  assign stOp_lane[10].cntl__stOp__strm0_source       = cntl__sdp__lane10_strm0_stOp_source      ;
  assign stOp_lane[10].cntl__stOp__strm0_destination  = cntl__sdp__lane10_strm0_stOp_destination ;
  assign stOp_lane[10].cntl__stOp__strm1_source       = cntl__sdp__lane10_strm1_stOp_source      ;
  assign stOp_lane[10].cntl__stOp__strm1_destination  = cntl__sdp__lane10_strm1_stOp_destination ;
  assign stOp_lane[10].cntl__stOp__strm0_enable       = cntl__sdp__lane10_strm0_stOp_enable      ;
  assign sdp__cntl__lane10_strm0_stOp_ready           = stOp_lane[10].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane10_strm0_stOp_complete        = stOp_lane[10].stOp__cntl__strm0_complete ;
  assign stOp_lane[10].cntl__stOp__strm1_enable       = cntl__sdp__lane10_strm1_stOp_enable      ;
  assign sdp__cntl__lane10_strm1_stOp_ready           = stOp_lane[10].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane10_strm1_stOp_complete        = stOp_lane[10].stOp__cntl__strm1_complete ;
  assign stOp_lane[11].cntl__stOp__operation    = cntl__sdp__lane11_stOp_operation   ;
  assign stOp_lane[11].cntl__stOp__strm0_source       = cntl__sdp__lane11_strm0_stOp_source      ;
  assign stOp_lane[11].cntl__stOp__strm0_destination  = cntl__sdp__lane11_strm0_stOp_destination ;
  assign stOp_lane[11].cntl__stOp__strm1_source       = cntl__sdp__lane11_strm1_stOp_source      ;
  assign stOp_lane[11].cntl__stOp__strm1_destination  = cntl__sdp__lane11_strm1_stOp_destination ;
  assign stOp_lane[11].cntl__stOp__strm0_enable       = cntl__sdp__lane11_strm0_stOp_enable      ;
  assign sdp__cntl__lane11_strm0_stOp_ready           = stOp_lane[11].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane11_strm0_stOp_complete        = stOp_lane[11].stOp__cntl__strm0_complete ;
  assign stOp_lane[11].cntl__stOp__strm1_enable       = cntl__sdp__lane11_strm1_stOp_enable      ;
  assign sdp__cntl__lane11_strm1_stOp_ready           = stOp_lane[11].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane11_strm1_stOp_complete        = stOp_lane[11].stOp__cntl__strm1_complete ;
  assign stOp_lane[12].cntl__stOp__operation    = cntl__sdp__lane12_stOp_operation   ;
  assign stOp_lane[12].cntl__stOp__strm0_source       = cntl__sdp__lane12_strm0_stOp_source      ;
  assign stOp_lane[12].cntl__stOp__strm0_destination  = cntl__sdp__lane12_strm0_stOp_destination ;
  assign stOp_lane[12].cntl__stOp__strm1_source       = cntl__sdp__lane12_strm1_stOp_source      ;
  assign stOp_lane[12].cntl__stOp__strm1_destination  = cntl__sdp__lane12_strm1_stOp_destination ;
  assign stOp_lane[12].cntl__stOp__strm0_enable       = cntl__sdp__lane12_strm0_stOp_enable      ;
  assign sdp__cntl__lane12_strm0_stOp_ready           = stOp_lane[12].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane12_strm0_stOp_complete        = stOp_lane[12].stOp__cntl__strm0_complete ;
  assign stOp_lane[12].cntl__stOp__strm1_enable       = cntl__sdp__lane12_strm1_stOp_enable      ;
  assign sdp__cntl__lane12_strm1_stOp_ready           = stOp_lane[12].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane12_strm1_stOp_complete        = stOp_lane[12].stOp__cntl__strm1_complete ;
  assign stOp_lane[13].cntl__stOp__operation    = cntl__sdp__lane13_stOp_operation   ;
  assign stOp_lane[13].cntl__stOp__strm0_source       = cntl__sdp__lane13_strm0_stOp_source      ;
  assign stOp_lane[13].cntl__stOp__strm0_destination  = cntl__sdp__lane13_strm0_stOp_destination ;
  assign stOp_lane[13].cntl__stOp__strm1_source       = cntl__sdp__lane13_strm1_stOp_source      ;
  assign stOp_lane[13].cntl__stOp__strm1_destination  = cntl__sdp__lane13_strm1_stOp_destination ;
  assign stOp_lane[13].cntl__stOp__strm0_enable       = cntl__sdp__lane13_strm0_stOp_enable      ;
  assign sdp__cntl__lane13_strm0_stOp_ready           = stOp_lane[13].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane13_strm0_stOp_complete        = stOp_lane[13].stOp__cntl__strm0_complete ;
  assign stOp_lane[13].cntl__stOp__strm1_enable       = cntl__sdp__lane13_strm1_stOp_enable      ;
  assign sdp__cntl__lane13_strm1_stOp_ready           = stOp_lane[13].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane13_strm1_stOp_complete        = stOp_lane[13].stOp__cntl__strm1_complete ;
  assign stOp_lane[14].cntl__stOp__operation    = cntl__sdp__lane14_stOp_operation   ;
  assign stOp_lane[14].cntl__stOp__strm0_source       = cntl__sdp__lane14_strm0_stOp_source      ;
  assign stOp_lane[14].cntl__stOp__strm0_destination  = cntl__sdp__lane14_strm0_stOp_destination ;
  assign stOp_lane[14].cntl__stOp__strm1_source       = cntl__sdp__lane14_strm1_stOp_source      ;
  assign stOp_lane[14].cntl__stOp__strm1_destination  = cntl__sdp__lane14_strm1_stOp_destination ;
  assign stOp_lane[14].cntl__stOp__strm0_enable       = cntl__sdp__lane14_strm0_stOp_enable      ;
  assign sdp__cntl__lane14_strm0_stOp_ready           = stOp_lane[14].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane14_strm0_stOp_complete        = stOp_lane[14].stOp__cntl__strm0_complete ;
  assign stOp_lane[14].cntl__stOp__strm1_enable       = cntl__sdp__lane14_strm1_stOp_enable      ;
  assign sdp__cntl__lane14_strm1_stOp_ready           = stOp_lane[14].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane14_strm1_stOp_complete        = stOp_lane[14].stOp__cntl__strm1_complete ;
  assign stOp_lane[15].cntl__stOp__operation    = cntl__sdp__lane15_stOp_operation   ;
  assign stOp_lane[15].cntl__stOp__strm0_source       = cntl__sdp__lane15_strm0_stOp_source      ;
  assign stOp_lane[15].cntl__stOp__strm0_destination  = cntl__sdp__lane15_strm0_stOp_destination ;
  assign stOp_lane[15].cntl__stOp__strm1_source       = cntl__sdp__lane15_strm1_stOp_source      ;
  assign stOp_lane[15].cntl__stOp__strm1_destination  = cntl__sdp__lane15_strm1_stOp_destination ;
  assign stOp_lane[15].cntl__stOp__strm0_enable       = cntl__sdp__lane15_strm0_stOp_enable      ;
  assign sdp__cntl__lane15_strm0_stOp_ready           = stOp_lane[15].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane15_strm0_stOp_complete        = stOp_lane[15].stOp__cntl__strm0_complete ;
  assign stOp_lane[15].cntl__stOp__strm1_enable       = cntl__sdp__lane15_strm1_stOp_enable      ;
  assign sdp__cntl__lane15_strm1_stOp_ready           = stOp_lane[15].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane15_strm1_stOp_complete        = stOp_lane[15].stOp__cntl__strm1_complete ;
  assign stOp_lane[16].cntl__stOp__operation    = cntl__sdp__lane16_stOp_operation   ;
  assign stOp_lane[16].cntl__stOp__strm0_source       = cntl__sdp__lane16_strm0_stOp_source      ;
  assign stOp_lane[16].cntl__stOp__strm0_destination  = cntl__sdp__lane16_strm0_stOp_destination ;
  assign stOp_lane[16].cntl__stOp__strm1_source       = cntl__sdp__lane16_strm1_stOp_source      ;
  assign stOp_lane[16].cntl__stOp__strm1_destination  = cntl__sdp__lane16_strm1_stOp_destination ;
  assign stOp_lane[16].cntl__stOp__strm0_enable       = cntl__sdp__lane16_strm0_stOp_enable      ;
  assign sdp__cntl__lane16_strm0_stOp_ready           = stOp_lane[16].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane16_strm0_stOp_complete        = stOp_lane[16].stOp__cntl__strm0_complete ;
  assign stOp_lane[16].cntl__stOp__strm1_enable       = cntl__sdp__lane16_strm1_stOp_enable      ;
  assign sdp__cntl__lane16_strm1_stOp_ready           = stOp_lane[16].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane16_strm1_stOp_complete        = stOp_lane[16].stOp__cntl__strm1_complete ;
  assign stOp_lane[17].cntl__stOp__operation    = cntl__sdp__lane17_stOp_operation   ;
  assign stOp_lane[17].cntl__stOp__strm0_source       = cntl__sdp__lane17_strm0_stOp_source      ;
  assign stOp_lane[17].cntl__stOp__strm0_destination  = cntl__sdp__lane17_strm0_stOp_destination ;
  assign stOp_lane[17].cntl__stOp__strm1_source       = cntl__sdp__lane17_strm1_stOp_source      ;
  assign stOp_lane[17].cntl__stOp__strm1_destination  = cntl__sdp__lane17_strm1_stOp_destination ;
  assign stOp_lane[17].cntl__stOp__strm0_enable       = cntl__sdp__lane17_strm0_stOp_enable      ;
  assign sdp__cntl__lane17_strm0_stOp_ready           = stOp_lane[17].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane17_strm0_stOp_complete        = stOp_lane[17].stOp__cntl__strm0_complete ;
  assign stOp_lane[17].cntl__stOp__strm1_enable       = cntl__sdp__lane17_strm1_stOp_enable      ;
  assign sdp__cntl__lane17_strm1_stOp_ready           = stOp_lane[17].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane17_strm1_stOp_complete        = stOp_lane[17].stOp__cntl__strm1_complete ;
  assign stOp_lane[18].cntl__stOp__operation    = cntl__sdp__lane18_stOp_operation   ;
  assign stOp_lane[18].cntl__stOp__strm0_source       = cntl__sdp__lane18_strm0_stOp_source      ;
  assign stOp_lane[18].cntl__stOp__strm0_destination  = cntl__sdp__lane18_strm0_stOp_destination ;
  assign stOp_lane[18].cntl__stOp__strm1_source       = cntl__sdp__lane18_strm1_stOp_source      ;
  assign stOp_lane[18].cntl__stOp__strm1_destination  = cntl__sdp__lane18_strm1_stOp_destination ;
  assign stOp_lane[18].cntl__stOp__strm0_enable       = cntl__sdp__lane18_strm0_stOp_enable      ;
  assign sdp__cntl__lane18_strm0_stOp_ready           = stOp_lane[18].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane18_strm0_stOp_complete        = stOp_lane[18].stOp__cntl__strm0_complete ;
  assign stOp_lane[18].cntl__stOp__strm1_enable       = cntl__sdp__lane18_strm1_stOp_enable      ;
  assign sdp__cntl__lane18_strm1_stOp_ready           = stOp_lane[18].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane18_strm1_stOp_complete        = stOp_lane[18].stOp__cntl__strm1_complete ;
  assign stOp_lane[19].cntl__stOp__operation    = cntl__sdp__lane19_stOp_operation   ;
  assign stOp_lane[19].cntl__stOp__strm0_source       = cntl__sdp__lane19_strm0_stOp_source      ;
  assign stOp_lane[19].cntl__stOp__strm0_destination  = cntl__sdp__lane19_strm0_stOp_destination ;
  assign stOp_lane[19].cntl__stOp__strm1_source       = cntl__sdp__lane19_strm1_stOp_source      ;
  assign stOp_lane[19].cntl__stOp__strm1_destination  = cntl__sdp__lane19_strm1_stOp_destination ;
  assign stOp_lane[19].cntl__stOp__strm0_enable       = cntl__sdp__lane19_strm0_stOp_enable      ;
  assign sdp__cntl__lane19_strm0_stOp_ready           = stOp_lane[19].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane19_strm0_stOp_complete        = stOp_lane[19].stOp__cntl__strm0_complete ;
  assign stOp_lane[19].cntl__stOp__strm1_enable       = cntl__sdp__lane19_strm1_stOp_enable      ;
  assign sdp__cntl__lane19_strm1_stOp_ready           = stOp_lane[19].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane19_strm1_stOp_complete        = stOp_lane[19].stOp__cntl__strm1_complete ;
  assign stOp_lane[20].cntl__stOp__operation    = cntl__sdp__lane20_stOp_operation   ;
  assign stOp_lane[20].cntl__stOp__strm0_source       = cntl__sdp__lane20_strm0_stOp_source      ;
  assign stOp_lane[20].cntl__stOp__strm0_destination  = cntl__sdp__lane20_strm0_stOp_destination ;
  assign stOp_lane[20].cntl__stOp__strm1_source       = cntl__sdp__lane20_strm1_stOp_source      ;
  assign stOp_lane[20].cntl__stOp__strm1_destination  = cntl__sdp__lane20_strm1_stOp_destination ;
  assign stOp_lane[20].cntl__stOp__strm0_enable       = cntl__sdp__lane20_strm0_stOp_enable      ;
  assign sdp__cntl__lane20_strm0_stOp_ready           = stOp_lane[20].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane20_strm0_stOp_complete        = stOp_lane[20].stOp__cntl__strm0_complete ;
  assign stOp_lane[20].cntl__stOp__strm1_enable       = cntl__sdp__lane20_strm1_stOp_enable      ;
  assign sdp__cntl__lane20_strm1_stOp_ready           = stOp_lane[20].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane20_strm1_stOp_complete        = stOp_lane[20].stOp__cntl__strm1_complete ;
  assign stOp_lane[21].cntl__stOp__operation    = cntl__sdp__lane21_stOp_operation   ;
  assign stOp_lane[21].cntl__stOp__strm0_source       = cntl__sdp__lane21_strm0_stOp_source      ;
  assign stOp_lane[21].cntl__stOp__strm0_destination  = cntl__sdp__lane21_strm0_stOp_destination ;
  assign stOp_lane[21].cntl__stOp__strm1_source       = cntl__sdp__lane21_strm1_stOp_source      ;
  assign stOp_lane[21].cntl__stOp__strm1_destination  = cntl__sdp__lane21_strm1_stOp_destination ;
  assign stOp_lane[21].cntl__stOp__strm0_enable       = cntl__sdp__lane21_strm0_stOp_enable      ;
  assign sdp__cntl__lane21_strm0_stOp_ready           = stOp_lane[21].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane21_strm0_stOp_complete        = stOp_lane[21].stOp__cntl__strm0_complete ;
  assign stOp_lane[21].cntl__stOp__strm1_enable       = cntl__sdp__lane21_strm1_stOp_enable      ;
  assign sdp__cntl__lane21_strm1_stOp_ready           = stOp_lane[21].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane21_strm1_stOp_complete        = stOp_lane[21].stOp__cntl__strm1_complete ;
  assign stOp_lane[22].cntl__stOp__operation    = cntl__sdp__lane22_stOp_operation   ;
  assign stOp_lane[22].cntl__stOp__strm0_source       = cntl__sdp__lane22_strm0_stOp_source      ;
  assign stOp_lane[22].cntl__stOp__strm0_destination  = cntl__sdp__lane22_strm0_stOp_destination ;
  assign stOp_lane[22].cntl__stOp__strm1_source       = cntl__sdp__lane22_strm1_stOp_source      ;
  assign stOp_lane[22].cntl__stOp__strm1_destination  = cntl__sdp__lane22_strm1_stOp_destination ;
  assign stOp_lane[22].cntl__stOp__strm0_enable       = cntl__sdp__lane22_strm0_stOp_enable      ;
  assign sdp__cntl__lane22_strm0_stOp_ready           = stOp_lane[22].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane22_strm0_stOp_complete        = stOp_lane[22].stOp__cntl__strm0_complete ;
  assign stOp_lane[22].cntl__stOp__strm1_enable       = cntl__sdp__lane22_strm1_stOp_enable      ;
  assign sdp__cntl__lane22_strm1_stOp_ready           = stOp_lane[22].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane22_strm1_stOp_complete        = stOp_lane[22].stOp__cntl__strm1_complete ;
  assign stOp_lane[23].cntl__stOp__operation    = cntl__sdp__lane23_stOp_operation   ;
  assign stOp_lane[23].cntl__stOp__strm0_source       = cntl__sdp__lane23_strm0_stOp_source      ;
  assign stOp_lane[23].cntl__stOp__strm0_destination  = cntl__sdp__lane23_strm0_stOp_destination ;
  assign stOp_lane[23].cntl__stOp__strm1_source       = cntl__sdp__lane23_strm1_stOp_source      ;
  assign stOp_lane[23].cntl__stOp__strm1_destination  = cntl__sdp__lane23_strm1_stOp_destination ;
  assign stOp_lane[23].cntl__stOp__strm0_enable       = cntl__sdp__lane23_strm0_stOp_enable      ;
  assign sdp__cntl__lane23_strm0_stOp_ready           = stOp_lane[23].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane23_strm0_stOp_complete        = stOp_lane[23].stOp__cntl__strm0_complete ;
  assign stOp_lane[23].cntl__stOp__strm1_enable       = cntl__sdp__lane23_strm1_stOp_enable      ;
  assign sdp__cntl__lane23_strm1_stOp_ready           = stOp_lane[23].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane23_strm1_stOp_complete        = stOp_lane[23].stOp__cntl__strm1_complete ;
  assign stOp_lane[24].cntl__stOp__operation    = cntl__sdp__lane24_stOp_operation   ;
  assign stOp_lane[24].cntl__stOp__strm0_source       = cntl__sdp__lane24_strm0_stOp_source      ;
  assign stOp_lane[24].cntl__stOp__strm0_destination  = cntl__sdp__lane24_strm0_stOp_destination ;
  assign stOp_lane[24].cntl__stOp__strm1_source       = cntl__sdp__lane24_strm1_stOp_source      ;
  assign stOp_lane[24].cntl__stOp__strm1_destination  = cntl__sdp__lane24_strm1_stOp_destination ;
  assign stOp_lane[24].cntl__stOp__strm0_enable       = cntl__sdp__lane24_strm0_stOp_enable      ;
  assign sdp__cntl__lane24_strm0_stOp_ready           = stOp_lane[24].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane24_strm0_stOp_complete        = stOp_lane[24].stOp__cntl__strm0_complete ;
  assign stOp_lane[24].cntl__stOp__strm1_enable       = cntl__sdp__lane24_strm1_stOp_enable      ;
  assign sdp__cntl__lane24_strm1_stOp_ready           = stOp_lane[24].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane24_strm1_stOp_complete        = stOp_lane[24].stOp__cntl__strm1_complete ;
  assign stOp_lane[25].cntl__stOp__operation    = cntl__sdp__lane25_stOp_operation   ;
  assign stOp_lane[25].cntl__stOp__strm0_source       = cntl__sdp__lane25_strm0_stOp_source      ;
  assign stOp_lane[25].cntl__stOp__strm0_destination  = cntl__sdp__lane25_strm0_stOp_destination ;
  assign stOp_lane[25].cntl__stOp__strm1_source       = cntl__sdp__lane25_strm1_stOp_source      ;
  assign stOp_lane[25].cntl__stOp__strm1_destination  = cntl__sdp__lane25_strm1_stOp_destination ;
  assign stOp_lane[25].cntl__stOp__strm0_enable       = cntl__sdp__lane25_strm0_stOp_enable      ;
  assign sdp__cntl__lane25_strm0_stOp_ready           = stOp_lane[25].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane25_strm0_stOp_complete        = stOp_lane[25].stOp__cntl__strm0_complete ;
  assign stOp_lane[25].cntl__stOp__strm1_enable       = cntl__sdp__lane25_strm1_stOp_enable      ;
  assign sdp__cntl__lane25_strm1_stOp_ready           = stOp_lane[25].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane25_strm1_stOp_complete        = stOp_lane[25].stOp__cntl__strm1_complete ;
  assign stOp_lane[26].cntl__stOp__operation    = cntl__sdp__lane26_stOp_operation   ;
  assign stOp_lane[26].cntl__stOp__strm0_source       = cntl__sdp__lane26_strm0_stOp_source      ;
  assign stOp_lane[26].cntl__stOp__strm0_destination  = cntl__sdp__lane26_strm0_stOp_destination ;
  assign stOp_lane[26].cntl__stOp__strm1_source       = cntl__sdp__lane26_strm1_stOp_source      ;
  assign stOp_lane[26].cntl__stOp__strm1_destination  = cntl__sdp__lane26_strm1_stOp_destination ;
  assign stOp_lane[26].cntl__stOp__strm0_enable       = cntl__sdp__lane26_strm0_stOp_enable      ;
  assign sdp__cntl__lane26_strm0_stOp_ready           = stOp_lane[26].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane26_strm0_stOp_complete        = stOp_lane[26].stOp__cntl__strm0_complete ;
  assign stOp_lane[26].cntl__stOp__strm1_enable       = cntl__sdp__lane26_strm1_stOp_enable      ;
  assign sdp__cntl__lane26_strm1_stOp_ready           = stOp_lane[26].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane26_strm1_stOp_complete        = stOp_lane[26].stOp__cntl__strm1_complete ;
  assign stOp_lane[27].cntl__stOp__operation    = cntl__sdp__lane27_stOp_operation   ;
  assign stOp_lane[27].cntl__stOp__strm0_source       = cntl__sdp__lane27_strm0_stOp_source      ;
  assign stOp_lane[27].cntl__stOp__strm0_destination  = cntl__sdp__lane27_strm0_stOp_destination ;
  assign stOp_lane[27].cntl__stOp__strm1_source       = cntl__sdp__lane27_strm1_stOp_source      ;
  assign stOp_lane[27].cntl__stOp__strm1_destination  = cntl__sdp__lane27_strm1_stOp_destination ;
  assign stOp_lane[27].cntl__stOp__strm0_enable       = cntl__sdp__lane27_strm0_stOp_enable      ;
  assign sdp__cntl__lane27_strm0_stOp_ready           = stOp_lane[27].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane27_strm0_stOp_complete        = stOp_lane[27].stOp__cntl__strm0_complete ;
  assign stOp_lane[27].cntl__stOp__strm1_enable       = cntl__sdp__lane27_strm1_stOp_enable      ;
  assign sdp__cntl__lane27_strm1_stOp_ready           = stOp_lane[27].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane27_strm1_stOp_complete        = stOp_lane[27].stOp__cntl__strm1_complete ;
  assign stOp_lane[28].cntl__stOp__operation    = cntl__sdp__lane28_stOp_operation   ;
  assign stOp_lane[28].cntl__stOp__strm0_source       = cntl__sdp__lane28_strm0_stOp_source      ;
  assign stOp_lane[28].cntl__stOp__strm0_destination  = cntl__sdp__lane28_strm0_stOp_destination ;
  assign stOp_lane[28].cntl__stOp__strm1_source       = cntl__sdp__lane28_strm1_stOp_source      ;
  assign stOp_lane[28].cntl__stOp__strm1_destination  = cntl__sdp__lane28_strm1_stOp_destination ;
  assign stOp_lane[28].cntl__stOp__strm0_enable       = cntl__sdp__lane28_strm0_stOp_enable      ;
  assign sdp__cntl__lane28_strm0_stOp_ready           = stOp_lane[28].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane28_strm0_stOp_complete        = stOp_lane[28].stOp__cntl__strm0_complete ;
  assign stOp_lane[28].cntl__stOp__strm1_enable       = cntl__sdp__lane28_strm1_stOp_enable      ;
  assign sdp__cntl__lane28_strm1_stOp_ready           = stOp_lane[28].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane28_strm1_stOp_complete        = stOp_lane[28].stOp__cntl__strm1_complete ;
  assign stOp_lane[29].cntl__stOp__operation    = cntl__sdp__lane29_stOp_operation   ;
  assign stOp_lane[29].cntl__stOp__strm0_source       = cntl__sdp__lane29_strm0_stOp_source      ;
  assign stOp_lane[29].cntl__stOp__strm0_destination  = cntl__sdp__lane29_strm0_stOp_destination ;
  assign stOp_lane[29].cntl__stOp__strm1_source       = cntl__sdp__lane29_strm1_stOp_source      ;
  assign stOp_lane[29].cntl__stOp__strm1_destination  = cntl__sdp__lane29_strm1_stOp_destination ;
  assign stOp_lane[29].cntl__stOp__strm0_enable       = cntl__sdp__lane29_strm0_stOp_enable      ;
  assign sdp__cntl__lane29_strm0_stOp_ready           = stOp_lane[29].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane29_strm0_stOp_complete        = stOp_lane[29].stOp__cntl__strm0_complete ;
  assign stOp_lane[29].cntl__stOp__strm1_enable       = cntl__sdp__lane29_strm1_stOp_enable      ;
  assign sdp__cntl__lane29_strm1_stOp_ready           = stOp_lane[29].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane29_strm1_stOp_complete        = stOp_lane[29].stOp__cntl__strm1_complete ;
  assign stOp_lane[30].cntl__stOp__operation    = cntl__sdp__lane30_stOp_operation   ;
  assign stOp_lane[30].cntl__stOp__strm0_source       = cntl__sdp__lane30_strm0_stOp_source      ;
  assign stOp_lane[30].cntl__stOp__strm0_destination  = cntl__sdp__lane30_strm0_stOp_destination ;
  assign stOp_lane[30].cntl__stOp__strm1_source       = cntl__sdp__lane30_strm1_stOp_source      ;
  assign stOp_lane[30].cntl__stOp__strm1_destination  = cntl__sdp__lane30_strm1_stOp_destination ;
  assign stOp_lane[30].cntl__stOp__strm0_enable       = cntl__sdp__lane30_strm0_stOp_enable      ;
  assign sdp__cntl__lane30_strm0_stOp_ready           = stOp_lane[30].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane30_strm0_stOp_complete        = stOp_lane[30].stOp__cntl__strm0_complete ;
  assign stOp_lane[30].cntl__stOp__strm1_enable       = cntl__sdp__lane30_strm1_stOp_enable      ;
  assign sdp__cntl__lane30_strm1_stOp_ready           = stOp_lane[30].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane30_strm1_stOp_complete        = stOp_lane[30].stOp__cntl__strm1_complete ;
  assign stOp_lane[31].cntl__stOp__operation    = cntl__sdp__lane31_stOp_operation   ;
  assign stOp_lane[31].cntl__stOp__strm0_source       = cntl__sdp__lane31_strm0_stOp_source      ;
  assign stOp_lane[31].cntl__stOp__strm0_destination  = cntl__sdp__lane31_strm0_stOp_destination ;
  assign stOp_lane[31].cntl__stOp__strm1_source       = cntl__sdp__lane31_strm1_stOp_source      ;
  assign stOp_lane[31].cntl__stOp__strm1_destination  = cntl__sdp__lane31_strm1_stOp_destination ;
  assign stOp_lane[31].cntl__stOp__strm0_enable       = cntl__sdp__lane31_strm0_stOp_enable      ;
  assign sdp__cntl__lane31_strm0_stOp_ready           = stOp_lane[31].stOp__cntl__strm0_ready    ;
  assign sdp__cntl__lane31_strm0_stOp_complete        = stOp_lane[31].stOp__cntl__strm0_complete ;
  assign stOp_lane[31].cntl__stOp__strm1_enable       = cntl__sdp__lane31_strm1_stOp_enable      ;
  assign sdp__cntl__lane31_strm1_stOp_ready           = stOp_lane[31].stOp__cntl__strm1_ready    ;
  assign sdp__cntl__lane31_strm1_stOp_complete        = stOp_lane[31].stOp__cntl__strm1_complete ;
