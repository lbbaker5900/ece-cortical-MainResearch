
            begin
              @(final_operation[0][0]) ;
            end
            begin
              @(final_operation[0][1]) ;
            end
            begin
              @(final_operation[0][2]) ;
            end
            begin
              @(final_operation[0][3]) ;
            end
            begin
              @(final_operation[0][4]) ;
            end
            begin
              @(final_operation[0][5]) ;
            end
            begin
              @(final_operation[0][6]) ;
            end
            begin
              @(final_operation[0][7]) ;
            end
            begin
              @(final_operation[0][8]) ;
            end
            begin
              @(final_operation[0][9]) ;
            end
            begin
              @(final_operation[0][10]) ;
            end
            begin
              @(final_operation[0][11]) ;
            end
            begin
              @(final_operation[0][12]) ;
            end
            begin
              @(final_operation[0][13]) ;
            end
            begin
              @(final_operation[0][14]) ;
            end
            begin
              @(final_operation[0][15]) ;
            end
            begin
              @(final_operation[0][16]) ;
            end
            begin
              @(final_operation[0][17]) ;
            end
            begin
              @(final_operation[0][18]) ;
            end
            begin
              @(final_operation[0][19]) ;
            end
            begin
              @(final_operation[0][20]) ;
            end
            begin
              @(final_operation[0][21]) ;
            end
            begin
              @(final_operation[0][22]) ;
            end
            begin
              @(final_operation[0][23]) ;
            end
            begin
              @(final_operation[0][24]) ;
            end
            begin
              @(final_operation[0][25]) ;
            end
            begin
              @(final_operation[0][26]) ;
            end
            begin
              @(final_operation[0][27]) ;
            end
            begin
              @(final_operation[0][28]) ;
            end
            begin
              @(final_operation[0][29]) ;
            end
            begin
              @(final_operation[0][30]) ;
            end
            begin
              @(final_operation[0][31]) ;
            end

            begin
              @(final_operation[1][0]) ;
            end
            begin
              @(final_operation[1][1]) ;
            end
            begin
              @(final_operation[1][2]) ;
            end
            begin
              @(final_operation[1][3]) ;
            end
            begin
              @(final_operation[1][4]) ;
            end
            begin
              @(final_operation[1][5]) ;
            end
            begin
              @(final_operation[1][6]) ;
            end
            begin
              @(final_operation[1][7]) ;
            end
            begin
              @(final_operation[1][8]) ;
            end
            begin
              @(final_operation[1][9]) ;
            end
            begin
              @(final_operation[1][10]) ;
            end
            begin
              @(final_operation[1][11]) ;
            end
            begin
              @(final_operation[1][12]) ;
            end
            begin
              @(final_operation[1][13]) ;
            end
            begin
              @(final_operation[1][14]) ;
            end
            begin
              @(final_operation[1][15]) ;
            end
            begin
              @(final_operation[1][16]) ;
            end
            begin
              @(final_operation[1][17]) ;
            end
            begin
              @(final_operation[1][18]) ;
            end
            begin
              @(final_operation[1][19]) ;
            end
            begin
              @(final_operation[1][20]) ;
            end
            begin
              @(final_operation[1][21]) ;
            end
            begin
              @(final_operation[1][22]) ;
            end
            begin
              @(final_operation[1][23]) ;
            end
            begin
              @(final_operation[1][24]) ;
            end
            begin
              @(final_operation[1][25]) ;
            end
            begin
              @(final_operation[1][26]) ;
            end
            begin
              @(final_operation[1][27]) ;
            end
            begin
              @(final_operation[1][28]) ;
            end
            begin
              @(final_operation[1][29]) ;
            end
            begin
              @(final_operation[1][30]) ;
            end
            begin
              @(final_operation[1][31]) ;
            end

            begin
              @(final_operation[2][0]) ;
            end
            begin
              @(final_operation[2][1]) ;
            end
            begin
              @(final_operation[2][2]) ;
            end
            begin
              @(final_operation[2][3]) ;
            end
            begin
              @(final_operation[2][4]) ;
            end
            begin
              @(final_operation[2][5]) ;
            end
            begin
              @(final_operation[2][6]) ;
            end
            begin
              @(final_operation[2][7]) ;
            end
            begin
              @(final_operation[2][8]) ;
            end
            begin
              @(final_operation[2][9]) ;
            end
            begin
              @(final_operation[2][10]) ;
            end
            begin
              @(final_operation[2][11]) ;
            end
            begin
              @(final_operation[2][12]) ;
            end
            begin
              @(final_operation[2][13]) ;
            end
            begin
              @(final_operation[2][14]) ;
            end
            begin
              @(final_operation[2][15]) ;
            end
            begin
              @(final_operation[2][16]) ;
            end
            begin
              @(final_operation[2][17]) ;
            end
            begin
              @(final_operation[2][18]) ;
            end
            begin
              @(final_operation[2][19]) ;
            end
            begin
              @(final_operation[2][20]) ;
            end
            begin
              @(final_operation[2][21]) ;
            end
            begin
              @(final_operation[2][22]) ;
            end
            begin
              @(final_operation[2][23]) ;
            end
            begin
              @(final_operation[2][24]) ;
            end
            begin
              @(final_operation[2][25]) ;
            end
            begin
              @(final_operation[2][26]) ;
            end
            begin
              @(final_operation[2][27]) ;
            end
            begin
              @(final_operation[2][28]) ;
            end
            begin
              @(final_operation[2][29]) ;
            end
            begin
              @(final_operation[2][30]) ;
            end
            begin
              @(final_operation[2][31]) ;
            end

            begin
              @(final_operation[3][0]) ;
            end
            begin
              @(final_operation[3][1]) ;
            end
            begin
              @(final_operation[3][2]) ;
            end
            begin
              @(final_operation[3][3]) ;
            end
            begin
              @(final_operation[3][4]) ;
            end
            begin
              @(final_operation[3][5]) ;
            end
            begin
              @(final_operation[3][6]) ;
            end
            begin
              @(final_operation[3][7]) ;
            end
            begin
              @(final_operation[3][8]) ;
            end
            begin
              @(final_operation[3][9]) ;
            end
            begin
              @(final_operation[3][10]) ;
            end
            begin
              @(final_operation[3][11]) ;
            end
            begin
              @(final_operation[3][12]) ;
            end
            begin
              @(final_operation[3][13]) ;
            end
            begin
              @(final_operation[3][14]) ;
            end
            begin
              @(final_operation[3][15]) ;
            end
            begin
              @(final_operation[3][16]) ;
            end
            begin
              @(final_operation[3][17]) ;
            end
            begin
              @(final_operation[3][18]) ;
            end
            begin
              @(final_operation[3][19]) ;
            end
            begin
              @(final_operation[3][20]) ;
            end
            begin
              @(final_operation[3][21]) ;
            end
            begin
              @(final_operation[3][22]) ;
            end
            begin
              @(final_operation[3][23]) ;
            end
            begin
              @(final_operation[3][24]) ;
            end
            begin
              @(final_operation[3][25]) ;
            end
            begin
              @(final_operation[3][26]) ;
            end
            begin
              @(final_operation[3][27]) ;
            end
            begin
              @(final_operation[3][28]) ;
            end
            begin
              @(final_operation[3][29]) ;
            end
            begin
              @(final_operation[3][30]) ;
            end
            begin
              @(final_operation[3][31]) ;
            end

            begin
              @(final_operation[4][0]) ;
            end
            begin
              @(final_operation[4][1]) ;
            end
            begin
              @(final_operation[4][2]) ;
            end
            begin
              @(final_operation[4][3]) ;
            end
            begin
              @(final_operation[4][4]) ;
            end
            begin
              @(final_operation[4][5]) ;
            end
            begin
              @(final_operation[4][6]) ;
            end
            begin
              @(final_operation[4][7]) ;
            end
            begin
              @(final_operation[4][8]) ;
            end
            begin
              @(final_operation[4][9]) ;
            end
            begin
              @(final_operation[4][10]) ;
            end
            begin
              @(final_operation[4][11]) ;
            end
            begin
              @(final_operation[4][12]) ;
            end
            begin
              @(final_operation[4][13]) ;
            end
            begin
              @(final_operation[4][14]) ;
            end
            begin
              @(final_operation[4][15]) ;
            end
            begin
              @(final_operation[4][16]) ;
            end
            begin
              @(final_operation[4][17]) ;
            end
            begin
              @(final_operation[4][18]) ;
            end
            begin
              @(final_operation[4][19]) ;
            end
            begin
              @(final_operation[4][20]) ;
            end
            begin
              @(final_operation[4][21]) ;
            end
            begin
              @(final_operation[4][22]) ;
            end
            begin
              @(final_operation[4][23]) ;
            end
            begin
              @(final_operation[4][24]) ;
            end
            begin
              @(final_operation[4][25]) ;
            end
            begin
              @(final_operation[4][26]) ;
            end
            begin
              @(final_operation[4][27]) ;
            end
            begin
              @(final_operation[4][28]) ;
            end
            begin
              @(final_operation[4][29]) ;
            end
            begin
              @(final_operation[4][30]) ;
            end
            begin
              @(final_operation[4][31]) ;
            end

            begin
              @(final_operation[5][0]) ;
            end
            begin
              @(final_operation[5][1]) ;
            end
            begin
              @(final_operation[5][2]) ;
            end
            begin
              @(final_operation[5][3]) ;
            end
            begin
              @(final_operation[5][4]) ;
            end
            begin
              @(final_operation[5][5]) ;
            end
            begin
              @(final_operation[5][6]) ;
            end
            begin
              @(final_operation[5][7]) ;
            end
            begin
              @(final_operation[5][8]) ;
            end
            begin
              @(final_operation[5][9]) ;
            end
            begin
              @(final_operation[5][10]) ;
            end
            begin
              @(final_operation[5][11]) ;
            end
            begin
              @(final_operation[5][12]) ;
            end
            begin
              @(final_operation[5][13]) ;
            end
            begin
              @(final_operation[5][14]) ;
            end
            begin
              @(final_operation[5][15]) ;
            end
            begin
              @(final_operation[5][16]) ;
            end
            begin
              @(final_operation[5][17]) ;
            end
            begin
              @(final_operation[5][18]) ;
            end
            begin
              @(final_operation[5][19]) ;
            end
            begin
              @(final_operation[5][20]) ;
            end
            begin
              @(final_operation[5][21]) ;
            end
            begin
              @(final_operation[5][22]) ;
            end
            begin
              @(final_operation[5][23]) ;
            end
            begin
              @(final_operation[5][24]) ;
            end
            begin
              @(final_operation[5][25]) ;
            end
            begin
              @(final_operation[5][26]) ;
            end
            begin
              @(final_operation[5][27]) ;
            end
            begin
              @(final_operation[5][28]) ;
            end
            begin
              @(final_operation[5][29]) ;
            end
            begin
              @(final_operation[5][30]) ;
            end
            begin
              @(final_operation[5][31]) ;
            end

            begin
              @(final_operation[6][0]) ;
            end
            begin
              @(final_operation[6][1]) ;
            end
            begin
              @(final_operation[6][2]) ;
            end
            begin
              @(final_operation[6][3]) ;
            end
            begin
              @(final_operation[6][4]) ;
            end
            begin
              @(final_operation[6][5]) ;
            end
            begin
              @(final_operation[6][6]) ;
            end
            begin
              @(final_operation[6][7]) ;
            end
            begin
              @(final_operation[6][8]) ;
            end
            begin
              @(final_operation[6][9]) ;
            end
            begin
              @(final_operation[6][10]) ;
            end
            begin
              @(final_operation[6][11]) ;
            end
            begin
              @(final_operation[6][12]) ;
            end
            begin
              @(final_operation[6][13]) ;
            end
            begin
              @(final_operation[6][14]) ;
            end
            begin
              @(final_operation[6][15]) ;
            end
            begin
              @(final_operation[6][16]) ;
            end
            begin
              @(final_operation[6][17]) ;
            end
            begin
              @(final_operation[6][18]) ;
            end
            begin
              @(final_operation[6][19]) ;
            end
            begin
              @(final_operation[6][20]) ;
            end
            begin
              @(final_operation[6][21]) ;
            end
            begin
              @(final_operation[6][22]) ;
            end
            begin
              @(final_operation[6][23]) ;
            end
            begin
              @(final_operation[6][24]) ;
            end
            begin
              @(final_operation[6][25]) ;
            end
            begin
              @(final_operation[6][26]) ;
            end
            begin
              @(final_operation[6][27]) ;
            end
            begin
              @(final_operation[6][28]) ;
            end
            begin
              @(final_operation[6][29]) ;
            end
            begin
              @(final_operation[6][30]) ;
            end
            begin
              @(final_operation[6][31]) ;
            end

            begin
              @(final_operation[7][0]) ;
            end
            begin
              @(final_operation[7][1]) ;
            end
            begin
              @(final_operation[7][2]) ;
            end
            begin
              @(final_operation[7][3]) ;
            end
            begin
              @(final_operation[7][4]) ;
            end
            begin
              @(final_operation[7][5]) ;
            end
            begin
              @(final_operation[7][6]) ;
            end
            begin
              @(final_operation[7][7]) ;
            end
            begin
              @(final_operation[7][8]) ;
            end
            begin
              @(final_operation[7][9]) ;
            end
            begin
              @(final_operation[7][10]) ;
            end
            begin
              @(final_operation[7][11]) ;
            end
            begin
              @(final_operation[7][12]) ;
            end
            begin
              @(final_operation[7][13]) ;
            end
            begin
              @(final_operation[7][14]) ;
            end
            begin
              @(final_operation[7][15]) ;
            end
            begin
              @(final_operation[7][16]) ;
            end
            begin
              @(final_operation[7][17]) ;
            end
            begin
              @(final_operation[7][18]) ;
            end
            begin
              @(final_operation[7][19]) ;
            end
            begin
              @(final_operation[7][20]) ;
            end
            begin
              @(final_operation[7][21]) ;
            end
            begin
              @(final_operation[7][22]) ;
            end
            begin
              @(final_operation[7][23]) ;
            end
            begin
              @(final_operation[7][24]) ;
            end
            begin
              @(final_operation[7][25]) ;
            end
            begin
              @(final_operation[7][26]) ;
            end
            begin
              @(final_operation[7][27]) ;
            end
            begin
              @(final_operation[7][28]) ;
            end
            begin
              @(final_operation[7][29]) ;
            end
            begin
              @(final_operation[7][30]) ;
            end
            begin
              @(final_operation[7][31]) ;
            end

            begin
              @(final_operation[8][0]) ;
            end
            begin
              @(final_operation[8][1]) ;
            end
            begin
              @(final_operation[8][2]) ;
            end
            begin
              @(final_operation[8][3]) ;
            end
            begin
              @(final_operation[8][4]) ;
            end
            begin
              @(final_operation[8][5]) ;
            end
            begin
              @(final_operation[8][6]) ;
            end
            begin
              @(final_operation[8][7]) ;
            end
            begin
              @(final_operation[8][8]) ;
            end
            begin
              @(final_operation[8][9]) ;
            end
            begin
              @(final_operation[8][10]) ;
            end
            begin
              @(final_operation[8][11]) ;
            end
            begin
              @(final_operation[8][12]) ;
            end
            begin
              @(final_operation[8][13]) ;
            end
            begin
              @(final_operation[8][14]) ;
            end
            begin
              @(final_operation[8][15]) ;
            end
            begin
              @(final_operation[8][16]) ;
            end
            begin
              @(final_operation[8][17]) ;
            end
            begin
              @(final_operation[8][18]) ;
            end
            begin
              @(final_operation[8][19]) ;
            end
            begin
              @(final_operation[8][20]) ;
            end
            begin
              @(final_operation[8][21]) ;
            end
            begin
              @(final_operation[8][22]) ;
            end
            begin
              @(final_operation[8][23]) ;
            end
            begin
              @(final_operation[8][24]) ;
            end
            begin
              @(final_operation[8][25]) ;
            end
            begin
              @(final_operation[8][26]) ;
            end
            begin
              @(final_operation[8][27]) ;
            end
            begin
              @(final_operation[8][28]) ;
            end
            begin
              @(final_operation[8][29]) ;
            end
            begin
              @(final_operation[8][30]) ;
            end
            begin
              @(final_operation[8][31]) ;
            end

            begin
              @(final_operation[9][0]) ;
            end
            begin
              @(final_operation[9][1]) ;
            end
            begin
              @(final_operation[9][2]) ;
            end
            begin
              @(final_operation[9][3]) ;
            end
            begin
              @(final_operation[9][4]) ;
            end
            begin
              @(final_operation[9][5]) ;
            end
            begin
              @(final_operation[9][6]) ;
            end
            begin
              @(final_operation[9][7]) ;
            end
            begin
              @(final_operation[9][8]) ;
            end
            begin
              @(final_operation[9][9]) ;
            end
            begin
              @(final_operation[9][10]) ;
            end
            begin
              @(final_operation[9][11]) ;
            end
            begin
              @(final_operation[9][12]) ;
            end
            begin
              @(final_operation[9][13]) ;
            end
            begin
              @(final_operation[9][14]) ;
            end
            begin
              @(final_operation[9][15]) ;
            end
            begin
              @(final_operation[9][16]) ;
            end
            begin
              @(final_operation[9][17]) ;
            end
            begin
              @(final_operation[9][18]) ;
            end
            begin
              @(final_operation[9][19]) ;
            end
            begin
              @(final_operation[9][20]) ;
            end
            begin
              @(final_operation[9][21]) ;
            end
            begin
              @(final_operation[9][22]) ;
            end
            begin
              @(final_operation[9][23]) ;
            end
            begin
              @(final_operation[9][24]) ;
            end
            begin
              @(final_operation[9][25]) ;
            end
            begin
              @(final_operation[9][26]) ;
            end
            begin
              @(final_operation[9][27]) ;
            end
            begin
              @(final_operation[9][28]) ;
            end
            begin
              @(final_operation[9][29]) ;
            end
            begin
              @(final_operation[9][30]) ;
            end
            begin
              @(final_operation[9][31]) ;
            end

            begin
              @(final_operation[10][0]) ;
            end
            begin
              @(final_operation[10][1]) ;
            end
            begin
              @(final_operation[10][2]) ;
            end
            begin
              @(final_operation[10][3]) ;
            end
            begin
              @(final_operation[10][4]) ;
            end
            begin
              @(final_operation[10][5]) ;
            end
            begin
              @(final_operation[10][6]) ;
            end
            begin
              @(final_operation[10][7]) ;
            end
            begin
              @(final_operation[10][8]) ;
            end
            begin
              @(final_operation[10][9]) ;
            end
            begin
              @(final_operation[10][10]) ;
            end
            begin
              @(final_operation[10][11]) ;
            end
            begin
              @(final_operation[10][12]) ;
            end
            begin
              @(final_operation[10][13]) ;
            end
            begin
              @(final_operation[10][14]) ;
            end
            begin
              @(final_operation[10][15]) ;
            end
            begin
              @(final_operation[10][16]) ;
            end
            begin
              @(final_operation[10][17]) ;
            end
            begin
              @(final_operation[10][18]) ;
            end
            begin
              @(final_operation[10][19]) ;
            end
            begin
              @(final_operation[10][20]) ;
            end
            begin
              @(final_operation[10][21]) ;
            end
            begin
              @(final_operation[10][22]) ;
            end
            begin
              @(final_operation[10][23]) ;
            end
            begin
              @(final_operation[10][24]) ;
            end
            begin
              @(final_operation[10][25]) ;
            end
            begin
              @(final_operation[10][26]) ;
            end
            begin
              @(final_operation[10][27]) ;
            end
            begin
              @(final_operation[10][28]) ;
            end
            begin
              @(final_operation[10][29]) ;
            end
            begin
              @(final_operation[10][30]) ;
            end
            begin
              @(final_operation[10][31]) ;
            end

            begin
              @(final_operation[11][0]) ;
            end
            begin
              @(final_operation[11][1]) ;
            end
            begin
              @(final_operation[11][2]) ;
            end
            begin
              @(final_operation[11][3]) ;
            end
            begin
              @(final_operation[11][4]) ;
            end
            begin
              @(final_operation[11][5]) ;
            end
            begin
              @(final_operation[11][6]) ;
            end
            begin
              @(final_operation[11][7]) ;
            end
            begin
              @(final_operation[11][8]) ;
            end
            begin
              @(final_operation[11][9]) ;
            end
            begin
              @(final_operation[11][10]) ;
            end
            begin
              @(final_operation[11][11]) ;
            end
            begin
              @(final_operation[11][12]) ;
            end
            begin
              @(final_operation[11][13]) ;
            end
            begin
              @(final_operation[11][14]) ;
            end
            begin
              @(final_operation[11][15]) ;
            end
            begin
              @(final_operation[11][16]) ;
            end
            begin
              @(final_operation[11][17]) ;
            end
            begin
              @(final_operation[11][18]) ;
            end
            begin
              @(final_operation[11][19]) ;
            end
            begin
              @(final_operation[11][20]) ;
            end
            begin
              @(final_operation[11][21]) ;
            end
            begin
              @(final_operation[11][22]) ;
            end
            begin
              @(final_operation[11][23]) ;
            end
            begin
              @(final_operation[11][24]) ;
            end
            begin
              @(final_operation[11][25]) ;
            end
            begin
              @(final_operation[11][26]) ;
            end
            begin
              @(final_operation[11][27]) ;
            end
            begin
              @(final_operation[11][28]) ;
            end
            begin
              @(final_operation[11][29]) ;
            end
            begin
              @(final_operation[11][30]) ;
            end
            begin
              @(final_operation[11][31]) ;
            end

            begin
              @(final_operation[12][0]) ;
            end
            begin
              @(final_operation[12][1]) ;
            end
            begin
              @(final_operation[12][2]) ;
            end
            begin
              @(final_operation[12][3]) ;
            end
            begin
              @(final_operation[12][4]) ;
            end
            begin
              @(final_operation[12][5]) ;
            end
            begin
              @(final_operation[12][6]) ;
            end
            begin
              @(final_operation[12][7]) ;
            end
            begin
              @(final_operation[12][8]) ;
            end
            begin
              @(final_operation[12][9]) ;
            end
            begin
              @(final_operation[12][10]) ;
            end
            begin
              @(final_operation[12][11]) ;
            end
            begin
              @(final_operation[12][12]) ;
            end
            begin
              @(final_operation[12][13]) ;
            end
            begin
              @(final_operation[12][14]) ;
            end
            begin
              @(final_operation[12][15]) ;
            end
            begin
              @(final_operation[12][16]) ;
            end
            begin
              @(final_operation[12][17]) ;
            end
            begin
              @(final_operation[12][18]) ;
            end
            begin
              @(final_operation[12][19]) ;
            end
            begin
              @(final_operation[12][20]) ;
            end
            begin
              @(final_operation[12][21]) ;
            end
            begin
              @(final_operation[12][22]) ;
            end
            begin
              @(final_operation[12][23]) ;
            end
            begin
              @(final_operation[12][24]) ;
            end
            begin
              @(final_operation[12][25]) ;
            end
            begin
              @(final_operation[12][26]) ;
            end
            begin
              @(final_operation[12][27]) ;
            end
            begin
              @(final_operation[12][28]) ;
            end
            begin
              @(final_operation[12][29]) ;
            end
            begin
              @(final_operation[12][30]) ;
            end
            begin
              @(final_operation[12][31]) ;
            end

            begin
              @(final_operation[13][0]) ;
            end
            begin
              @(final_operation[13][1]) ;
            end
            begin
              @(final_operation[13][2]) ;
            end
            begin
              @(final_operation[13][3]) ;
            end
            begin
              @(final_operation[13][4]) ;
            end
            begin
              @(final_operation[13][5]) ;
            end
            begin
              @(final_operation[13][6]) ;
            end
            begin
              @(final_operation[13][7]) ;
            end
            begin
              @(final_operation[13][8]) ;
            end
            begin
              @(final_operation[13][9]) ;
            end
            begin
              @(final_operation[13][10]) ;
            end
            begin
              @(final_operation[13][11]) ;
            end
            begin
              @(final_operation[13][12]) ;
            end
            begin
              @(final_operation[13][13]) ;
            end
            begin
              @(final_operation[13][14]) ;
            end
            begin
              @(final_operation[13][15]) ;
            end
            begin
              @(final_operation[13][16]) ;
            end
            begin
              @(final_operation[13][17]) ;
            end
            begin
              @(final_operation[13][18]) ;
            end
            begin
              @(final_operation[13][19]) ;
            end
            begin
              @(final_operation[13][20]) ;
            end
            begin
              @(final_operation[13][21]) ;
            end
            begin
              @(final_operation[13][22]) ;
            end
            begin
              @(final_operation[13][23]) ;
            end
            begin
              @(final_operation[13][24]) ;
            end
            begin
              @(final_operation[13][25]) ;
            end
            begin
              @(final_operation[13][26]) ;
            end
            begin
              @(final_operation[13][27]) ;
            end
            begin
              @(final_operation[13][28]) ;
            end
            begin
              @(final_operation[13][29]) ;
            end
            begin
              @(final_operation[13][30]) ;
            end
            begin
              @(final_operation[13][31]) ;
            end

            begin
              @(final_operation[14][0]) ;
            end
            begin
              @(final_operation[14][1]) ;
            end
            begin
              @(final_operation[14][2]) ;
            end
            begin
              @(final_operation[14][3]) ;
            end
            begin
              @(final_operation[14][4]) ;
            end
            begin
              @(final_operation[14][5]) ;
            end
            begin
              @(final_operation[14][6]) ;
            end
            begin
              @(final_operation[14][7]) ;
            end
            begin
              @(final_operation[14][8]) ;
            end
            begin
              @(final_operation[14][9]) ;
            end
            begin
              @(final_operation[14][10]) ;
            end
            begin
              @(final_operation[14][11]) ;
            end
            begin
              @(final_operation[14][12]) ;
            end
            begin
              @(final_operation[14][13]) ;
            end
            begin
              @(final_operation[14][14]) ;
            end
            begin
              @(final_operation[14][15]) ;
            end
            begin
              @(final_operation[14][16]) ;
            end
            begin
              @(final_operation[14][17]) ;
            end
            begin
              @(final_operation[14][18]) ;
            end
            begin
              @(final_operation[14][19]) ;
            end
            begin
              @(final_operation[14][20]) ;
            end
            begin
              @(final_operation[14][21]) ;
            end
            begin
              @(final_operation[14][22]) ;
            end
            begin
              @(final_operation[14][23]) ;
            end
            begin
              @(final_operation[14][24]) ;
            end
            begin
              @(final_operation[14][25]) ;
            end
            begin
              @(final_operation[14][26]) ;
            end
            begin
              @(final_operation[14][27]) ;
            end
            begin
              @(final_operation[14][28]) ;
            end
            begin
              @(final_operation[14][29]) ;
            end
            begin
              @(final_operation[14][30]) ;
            end
            begin
              @(final_operation[14][31]) ;
            end

            begin
              @(final_operation[15][0]) ;
            end
            begin
              @(final_operation[15][1]) ;
            end
            begin
              @(final_operation[15][2]) ;
            end
            begin
              @(final_operation[15][3]) ;
            end
            begin
              @(final_operation[15][4]) ;
            end
            begin
              @(final_operation[15][5]) ;
            end
            begin
              @(final_operation[15][6]) ;
            end
            begin
              @(final_operation[15][7]) ;
            end
            begin
              @(final_operation[15][8]) ;
            end
            begin
              @(final_operation[15][9]) ;
            end
            begin
              @(final_operation[15][10]) ;
            end
            begin
              @(final_operation[15][11]) ;
            end
            begin
              @(final_operation[15][12]) ;
            end
            begin
              @(final_operation[15][13]) ;
            end
            begin
              @(final_operation[15][14]) ;
            end
            begin
              @(final_operation[15][15]) ;
            end
            begin
              @(final_operation[15][16]) ;
            end
            begin
              @(final_operation[15][17]) ;
            end
            begin
              @(final_operation[15][18]) ;
            end
            begin
              @(final_operation[15][19]) ;
            end
            begin
              @(final_operation[15][20]) ;
            end
            begin
              @(final_operation[15][21]) ;
            end
            begin
              @(final_operation[15][22]) ;
            end
            begin
              @(final_operation[15][23]) ;
            end
            begin
              @(final_operation[15][24]) ;
            end
            begin
              @(final_operation[15][25]) ;
            end
            begin
              @(final_operation[15][26]) ;
            end
            begin
              @(final_operation[15][27]) ;
            end
            begin
              @(final_operation[15][28]) ;
            end
            begin
              @(final_operation[15][29]) ;
            end
            begin
              @(final_operation[15][30]) ;
            end
            begin
              @(final_operation[15][31]) ;
            end

            begin
              @(final_operation[16][0]) ;
            end
            begin
              @(final_operation[16][1]) ;
            end
            begin
              @(final_operation[16][2]) ;
            end
            begin
              @(final_operation[16][3]) ;
            end
            begin
              @(final_operation[16][4]) ;
            end
            begin
              @(final_operation[16][5]) ;
            end
            begin
              @(final_operation[16][6]) ;
            end
            begin
              @(final_operation[16][7]) ;
            end
            begin
              @(final_operation[16][8]) ;
            end
            begin
              @(final_operation[16][9]) ;
            end
            begin
              @(final_operation[16][10]) ;
            end
            begin
              @(final_operation[16][11]) ;
            end
            begin
              @(final_operation[16][12]) ;
            end
            begin
              @(final_operation[16][13]) ;
            end
            begin
              @(final_operation[16][14]) ;
            end
            begin
              @(final_operation[16][15]) ;
            end
            begin
              @(final_operation[16][16]) ;
            end
            begin
              @(final_operation[16][17]) ;
            end
            begin
              @(final_operation[16][18]) ;
            end
            begin
              @(final_operation[16][19]) ;
            end
            begin
              @(final_operation[16][20]) ;
            end
            begin
              @(final_operation[16][21]) ;
            end
            begin
              @(final_operation[16][22]) ;
            end
            begin
              @(final_operation[16][23]) ;
            end
            begin
              @(final_operation[16][24]) ;
            end
            begin
              @(final_operation[16][25]) ;
            end
            begin
              @(final_operation[16][26]) ;
            end
            begin
              @(final_operation[16][27]) ;
            end
            begin
              @(final_operation[16][28]) ;
            end
            begin
              @(final_operation[16][29]) ;
            end
            begin
              @(final_operation[16][30]) ;
            end
            begin
              @(final_operation[16][31]) ;
            end

            begin
              @(final_operation[17][0]) ;
            end
            begin
              @(final_operation[17][1]) ;
            end
            begin
              @(final_operation[17][2]) ;
            end
            begin
              @(final_operation[17][3]) ;
            end
            begin
              @(final_operation[17][4]) ;
            end
            begin
              @(final_operation[17][5]) ;
            end
            begin
              @(final_operation[17][6]) ;
            end
            begin
              @(final_operation[17][7]) ;
            end
            begin
              @(final_operation[17][8]) ;
            end
            begin
              @(final_operation[17][9]) ;
            end
            begin
              @(final_operation[17][10]) ;
            end
            begin
              @(final_operation[17][11]) ;
            end
            begin
              @(final_operation[17][12]) ;
            end
            begin
              @(final_operation[17][13]) ;
            end
            begin
              @(final_operation[17][14]) ;
            end
            begin
              @(final_operation[17][15]) ;
            end
            begin
              @(final_operation[17][16]) ;
            end
            begin
              @(final_operation[17][17]) ;
            end
            begin
              @(final_operation[17][18]) ;
            end
            begin
              @(final_operation[17][19]) ;
            end
            begin
              @(final_operation[17][20]) ;
            end
            begin
              @(final_operation[17][21]) ;
            end
            begin
              @(final_operation[17][22]) ;
            end
            begin
              @(final_operation[17][23]) ;
            end
            begin
              @(final_operation[17][24]) ;
            end
            begin
              @(final_operation[17][25]) ;
            end
            begin
              @(final_operation[17][26]) ;
            end
            begin
              @(final_operation[17][27]) ;
            end
            begin
              @(final_operation[17][28]) ;
            end
            begin
              @(final_operation[17][29]) ;
            end
            begin
              @(final_operation[17][30]) ;
            end
            begin
              @(final_operation[17][31]) ;
            end

            begin
              @(final_operation[18][0]) ;
            end
            begin
              @(final_operation[18][1]) ;
            end
            begin
              @(final_operation[18][2]) ;
            end
            begin
              @(final_operation[18][3]) ;
            end
            begin
              @(final_operation[18][4]) ;
            end
            begin
              @(final_operation[18][5]) ;
            end
            begin
              @(final_operation[18][6]) ;
            end
            begin
              @(final_operation[18][7]) ;
            end
            begin
              @(final_operation[18][8]) ;
            end
            begin
              @(final_operation[18][9]) ;
            end
            begin
              @(final_operation[18][10]) ;
            end
            begin
              @(final_operation[18][11]) ;
            end
            begin
              @(final_operation[18][12]) ;
            end
            begin
              @(final_operation[18][13]) ;
            end
            begin
              @(final_operation[18][14]) ;
            end
            begin
              @(final_operation[18][15]) ;
            end
            begin
              @(final_operation[18][16]) ;
            end
            begin
              @(final_operation[18][17]) ;
            end
            begin
              @(final_operation[18][18]) ;
            end
            begin
              @(final_operation[18][19]) ;
            end
            begin
              @(final_operation[18][20]) ;
            end
            begin
              @(final_operation[18][21]) ;
            end
            begin
              @(final_operation[18][22]) ;
            end
            begin
              @(final_operation[18][23]) ;
            end
            begin
              @(final_operation[18][24]) ;
            end
            begin
              @(final_operation[18][25]) ;
            end
            begin
              @(final_operation[18][26]) ;
            end
            begin
              @(final_operation[18][27]) ;
            end
            begin
              @(final_operation[18][28]) ;
            end
            begin
              @(final_operation[18][29]) ;
            end
            begin
              @(final_operation[18][30]) ;
            end
            begin
              @(final_operation[18][31]) ;
            end

            begin
              @(final_operation[19][0]) ;
            end
            begin
              @(final_operation[19][1]) ;
            end
            begin
              @(final_operation[19][2]) ;
            end
            begin
              @(final_operation[19][3]) ;
            end
            begin
              @(final_operation[19][4]) ;
            end
            begin
              @(final_operation[19][5]) ;
            end
            begin
              @(final_operation[19][6]) ;
            end
            begin
              @(final_operation[19][7]) ;
            end
            begin
              @(final_operation[19][8]) ;
            end
            begin
              @(final_operation[19][9]) ;
            end
            begin
              @(final_operation[19][10]) ;
            end
            begin
              @(final_operation[19][11]) ;
            end
            begin
              @(final_operation[19][12]) ;
            end
            begin
              @(final_operation[19][13]) ;
            end
            begin
              @(final_operation[19][14]) ;
            end
            begin
              @(final_operation[19][15]) ;
            end
            begin
              @(final_operation[19][16]) ;
            end
            begin
              @(final_operation[19][17]) ;
            end
            begin
              @(final_operation[19][18]) ;
            end
            begin
              @(final_operation[19][19]) ;
            end
            begin
              @(final_operation[19][20]) ;
            end
            begin
              @(final_operation[19][21]) ;
            end
            begin
              @(final_operation[19][22]) ;
            end
            begin
              @(final_operation[19][23]) ;
            end
            begin
              @(final_operation[19][24]) ;
            end
            begin
              @(final_operation[19][25]) ;
            end
            begin
              @(final_operation[19][26]) ;
            end
            begin
              @(final_operation[19][27]) ;
            end
            begin
              @(final_operation[19][28]) ;
            end
            begin
              @(final_operation[19][29]) ;
            end
            begin
              @(final_operation[19][30]) ;
            end
            begin
              @(final_operation[19][31]) ;
            end

            begin
              @(final_operation[20][0]) ;
            end
            begin
              @(final_operation[20][1]) ;
            end
            begin
              @(final_operation[20][2]) ;
            end
            begin
              @(final_operation[20][3]) ;
            end
            begin
              @(final_operation[20][4]) ;
            end
            begin
              @(final_operation[20][5]) ;
            end
            begin
              @(final_operation[20][6]) ;
            end
            begin
              @(final_operation[20][7]) ;
            end
            begin
              @(final_operation[20][8]) ;
            end
            begin
              @(final_operation[20][9]) ;
            end
            begin
              @(final_operation[20][10]) ;
            end
            begin
              @(final_operation[20][11]) ;
            end
            begin
              @(final_operation[20][12]) ;
            end
            begin
              @(final_operation[20][13]) ;
            end
            begin
              @(final_operation[20][14]) ;
            end
            begin
              @(final_operation[20][15]) ;
            end
            begin
              @(final_operation[20][16]) ;
            end
            begin
              @(final_operation[20][17]) ;
            end
            begin
              @(final_operation[20][18]) ;
            end
            begin
              @(final_operation[20][19]) ;
            end
            begin
              @(final_operation[20][20]) ;
            end
            begin
              @(final_operation[20][21]) ;
            end
            begin
              @(final_operation[20][22]) ;
            end
            begin
              @(final_operation[20][23]) ;
            end
            begin
              @(final_operation[20][24]) ;
            end
            begin
              @(final_operation[20][25]) ;
            end
            begin
              @(final_operation[20][26]) ;
            end
            begin
              @(final_operation[20][27]) ;
            end
            begin
              @(final_operation[20][28]) ;
            end
            begin
              @(final_operation[20][29]) ;
            end
            begin
              @(final_operation[20][30]) ;
            end
            begin
              @(final_operation[20][31]) ;
            end

            begin
              @(final_operation[21][0]) ;
            end
            begin
              @(final_operation[21][1]) ;
            end
            begin
              @(final_operation[21][2]) ;
            end
            begin
              @(final_operation[21][3]) ;
            end
            begin
              @(final_operation[21][4]) ;
            end
            begin
              @(final_operation[21][5]) ;
            end
            begin
              @(final_operation[21][6]) ;
            end
            begin
              @(final_operation[21][7]) ;
            end
            begin
              @(final_operation[21][8]) ;
            end
            begin
              @(final_operation[21][9]) ;
            end
            begin
              @(final_operation[21][10]) ;
            end
            begin
              @(final_operation[21][11]) ;
            end
            begin
              @(final_operation[21][12]) ;
            end
            begin
              @(final_operation[21][13]) ;
            end
            begin
              @(final_operation[21][14]) ;
            end
            begin
              @(final_operation[21][15]) ;
            end
            begin
              @(final_operation[21][16]) ;
            end
            begin
              @(final_operation[21][17]) ;
            end
            begin
              @(final_operation[21][18]) ;
            end
            begin
              @(final_operation[21][19]) ;
            end
            begin
              @(final_operation[21][20]) ;
            end
            begin
              @(final_operation[21][21]) ;
            end
            begin
              @(final_operation[21][22]) ;
            end
            begin
              @(final_operation[21][23]) ;
            end
            begin
              @(final_operation[21][24]) ;
            end
            begin
              @(final_operation[21][25]) ;
            end
            begin
              @(final_operation[21][26]) ;
            end
            begin
              @(final_operation[21][27]) ;
            end
            begin
              @(final_operation[21][28]) ;
            end
            begin
              @(final_operation[21][29]) ;
            end
            begin
              @(final_operation[21][30]) ;
            end
            begin
              @(final_operation[21][31]) ;
            end

            begin
              @(final_operation[22][0]) ;
            end
            begin
              @(final_operation[22][1]) ;
            end
            begin
              @(final_operation[22][2]) ;
            end
            begin
              @(final_operation[22][3]) ;
            end
            begin
              @(final_operation[22][4]) ;
            end
            begin
              @(final_operation[22][5]) ;
            end
            begin
              @(final_operation[22][6]) ;
            end
            begin
              @(final_operation[22][7]) ;
            end
            begin
              @(final_operation[22][8]) ;
            end
            begin
              @(final_operation[22][9]) ;
            end
            begin
              @(final_operation[22][10]) ;
            end
            begin
              @(final_operation[22][11]) ;
            end
            begin
              @(final_operation[22][12]) ;
            end
            begin
              @(final_operation[22][13]) ;
            end
            begin
              @(final_operation[22][14]) ;
            end
            begin
              @(final_operation[22][15]) ;
            end
            begin
              @(final_operation[22][16]) ;
            end
            begin
              @(final_operation[22][17]) ;
            end
            begin
              @(final_operation[22][18]) ;
            end
            begin
              @(final_operation[22][19]) ;
            end
            begin
              @(final_operation[22][20]) ;
            end
            begin
              @(final_operation[22][21]) ;
            end
            begin
              @(final_operation[22][22]) ;
            end
            begin
              @(final_operation[22][23]) ;
            end
            begin
              @(final_operation[22][24]) ;
            end
            begin
              @(final_operation[22][25]) ;
            end
            begin
              @(final_operation[22][26]) ;
            end
            begin
              @(final_operation[22][27]) ;
            end
            begin
              @(final_operation[22][28]) ;
            end
            begin
              @(final_operation[22][29]) ;
            end
            begin
              @(final_operation[22][30]) ;
            end
            begin
              @(final_operation[22][31]) ;
            end

            begin
              @(final_operation[23][0]) ;
            end
            begin
              @(final_operation[23][1]) ;
            end
            begin
              @(final_operation[23][2]) ;
            end
            begin
              @(final_operation[23][3]) ;
            end
            begin
              @(final_operation[23][4]) ;
            end
            begin
              @(final_operation[23][5]) ;
            end
            begin
              @(final_operation[23][6]) ;
            end
            begin
              @(final_operation[23][7]) ;
            end
            begin
              @(final_operation[23][8]) ;
            end
            begin
              @(final_operation[23][9]) ;
            end
            begin
              @(final_operation[23][10]) ;
            end
            begin
              @(final_operation[23][11]) ;
            end
            begin
              @(final_operation[23][12]) ;
            end
            begin
              @(final_operation[23][13]) ;
            end
            begin
              @(final_operation[23][14]) ;
            end
            begin
              @(final_operation[23][15]) ;
            end
            begin
              @(final_operation[23][16]) ;
            end
            begin
              @(final_operation[23][17]) ;
            end
            begin
              @(final_operation[23][18]) ;
            end
            begin
              @(final_operation[23][19]) ;
            end
            begin
              @(final_operation[23][20]) ;
            end
            begin
              @(final_operation[23][21]) ;
            end
            begin
              @(final_operation[23][22]) ;
            end
            begin
              @(final_operation[23][23]) ;
            end
            begin
              @(final_operation[23][24]) ;
            end
            begin
              @(final_operation[23][25]) ;
            end
            begin
              @(final_operation[23][26]) ;
            end
            begin
              @(final_operation[23][27]) ;
            end
            begin
              @(final_operation[23][28]) ;
            end
            begin
              @(final_operation[23][29]) ;
            end
            begin
              @(final_operation[23][30]) ;
            end
            begin
              @(final_operation[23][31]) ;
            end

            begin
              @(final_operation[24][0]) ;
            end
            begin
              @(final_operation[24][1]) ;
            end
            begin
              @(final_operation[24][2]) ;
            end
            begin
              @(final_operation[24][3]) ;
            end
            begin
              @(final_operation[24][4]) ;
            end
            begin
              @(final_operation[24][5]) ;
            end
            begin
              @(final_operation[24][6]) ;
            end
            begin
              @(final_operation[24][7]) ;
            end
            begin
              @(final_operation[24][8]) ;
            end
            begin
              @(final_operation[24][9]) ;
            end
            begin
              @(final_operation[24][10]) ;
            end
            begin
              @(final_operation[24][11]) ;
            end
            begin
              @(final_operation[24][12]) ;
            end
            begin
              @(final_operation[24][13]) ;
            end
            begin
              @(final_operation[24][14]) ;
            end
            begin
              @(final_operation[24][15]) ;
            end
            begin
              @(final_operation[24][16]) ;
            end
            begin
              @(final_operation[24][17]) ;
            end
            begin
              @(final_operation[24][18]) ;
            end
            begin
              @(final_operation[24][19]) ;
            end
            begin
              @(final_operation[24][20]) ;
            end
            begin
              @(final_operation[24][21]) ;
            end
            begin
              @(final_operation[24][22]) ;
            end
            begin
              @(final_operation[24][23]) ;
            end
            begin
              @(final_operation[24][24]) ;
            end
            begin
              @(final_operation[24][25]) ;
            end
            begin
              @(final_operation[24][26]) ;
            end
            begin
              @(final_operation[24][27]) ;
            end
            begin
              @(final_operation[24][28]) ;
            end
            begin
              @(final_operation[24][29]) ;
            end
            begin
              @(final_operation[24][30]) ;
            end
            begin
              @(final_operation[24][31]) ;
            end

            begin
              @(final_operation[25][0]) ;
            end
            begin
              @(final_operation[25][1]) ;
            end
            begin
              @(final_operation[25][2]) ;
            end
            begin
              @(final_operation[25][3]) ;
            end
            begin
              @(final_operation[25][4]) ;
            end
            begin
              @(final_operation[25][5]) ;
            end
            begin
              @(final_operation[25][6]) ;
            end
            begin
              @(final_operation[25][7]) ;
            end
            begin
              @(final_operation[25][8]) ;
            end
            begin
              @(final_operation[25][9]) ;
            end
            begin
              @(final_operation[25][10]) ;
            end
            begin
              @(final_operation[25][11]) ;
            end
            begin
              @(final_operation[25][12]) ;
            end
            begin
              @(final_operation[25][13]) ;
            end
            begin
              @(final_operation[25][14]) ;
            end
            begin
              @(final_operation[25][15]) ;
            end
            begin
              @(final_operation[25][16]) ;
            end
            begin
              @(final_operation[25][17]) ;
            end
            begin
              @(final_operation[25][18]) ;
            end
            begin
              @(final_operation[25][19]) ;
            end
            begin
              @(final_operation[25][20]) ;
            end
            begin
              @(final_operation[25][21]) ;
            end
            begin
              @(final_operation[25][22]) ;
            end
            begin
              @(final_operation[25][23]) ;
            end
            begin
              @(final_operation[25][24]) ;
            end
            begin
              @(final_operation[25][25]) ;
            end
            begin
              @(final_operation[25][26]) ;
            end
            begin
              @(final_operation[25][27]) ;
            end
            begin
              @(final_operation[25][28]) ;
            end
            begin
              @(final_operation[25][29]) ;
            end
            begin
              @(final_operation[25][30]) ;
            end
            begin
              @(final_operation[25][31]) ;
            end

            begin
              @(final_operation[26][0]) ;
            end
            begin
              @(final_operation[26][1]) ;
            end
            begin
              @(final_operation[26][2]) ;
            end
            begin
              @(final_operation[26][3]) ;
            end
            begin
              @(final_operation[26][4]) ;
            end
            begin
              @(final_operation[26][5]) ;
            end
            begin
              @(final_operation[26][6]) ;
            end
            begin
              @(final_operation[26][7]) ;
            end
            begin
              @(final_operation[26][8]) ;
            end
            begin
              @(final_operation[26][9]) ;
            end
            begin
              @(final_operation[26][10]) ;
            end
            begin
              @(final_operation[26][11]) ;
            end
            begin
              @(final_operation[26][12]) ;
            end
            begin
              @(final_operation[26][13]) ;
            end
            begin
              @(final_operation[26][14]) ;
            end
            begin
              @(final_operation[26][15]) ;
            end
            begin
              @(final_operation[26][16]) ;
            end
            begin
              @(final_operation[26][17]) ;
            end
            begin
              @(final_operation[26][18]) ;
            end
            begin
              @(final_operation[26][19]) ;
            end
            begin
              @(final_operation[26][20]) ;
            end
            begin
              @(final_operation[26][21]) ;
            end
            begin
              @(final_operation[26][22]) ;
            end
            begin
              @(final_operation[26][23]) ;
            end
            begin
              @(final_operation[26][24]) ;
            end
            begin
              @(final_operation[26][25]) ;
            end
            begin
              @(final_operation[26][26]) ;
            end
            begin
              @(final_operation[26][27]) ;
            end
            begin
              @(final_operation[26][28]) ;
            end
            begin
              @(final_operation[26][29]) ;
            end
            begin
              @(final_operation[26][30]) ;
            end
            begin
              @(final_operation[26][31]) ;
            end

            begin
              @(final_operation[27][0]) ;
            end
            begin
              @(final_operation[27][1]) ;
            end
            begin
              @(final_operation[27][2]) ;
            end
            begin
              @(final_operation[27][3]) ;
            end
            begin
              @(final_operation[27][4]) ;
            end
            begin
              @(final_operation[27][5]) ;
            end
            begin
              @(final_operation[27][6]) ;
            end
            begin
              @(final_operation[27][7]) ;
            end
            begin
              @(final_operation[27][8]) ;
            end
            begin
              @(final_operation[27][9]) ;
            end
            begin
              @(final_operation[27][10]) ;
            end
            begin
              @(final_operation[27][11]) ;
            end
            begin
              @(final_operation[27][12]) ;
            end
            begin
              @(final_operation[27][13]) ;
            end
            begin
              @(final_operation[27][14]) ;
            end
            begin
              @(final_operation[27][15]) ;
            end
            begin
              @(final_operation[27][16]) ;
            end
            begin
              @(final_operation[27][17]) ;
            end
            begin
              @(final_operation[27][18]) ;
            end
            begin
              @(final_operation[27][19]) ;
            end
            begin
              @(final_operation[27][20]) ;
            end
            begin
              @(final_operation[27][21]) ;
            end
            begin
              @(final_operation[27][22]) ;
            end
            begin
              @(final_operation[27][23]) ;
            end
            begin
              @(final_operation[27][24]) ;
            end
            begin
              @(final_operation[27][25]) ;
            end
            begin
              @(final_operation[27][26]) ;
            end
            begin
              @(final_operation[27][27]) ;
            end
            begin
              @(final_operation[27][28]) ;
            end
            begin
              @(final_operation[27][29]) ;
            end
            begin
              @(final_operation[27][30]) ;
            end
            begin
              @(final_operation[27][31]) ;
            end

            begin
              @(final_operation[28][0]) ;
            end
            begin
              @(final_operation[28][1]) ;
            end
            begin
              @(final_operation[28][2]) ;
            end
            begin
              @(final_operation[28][3]) ;
            end
            begin
              @(final_operation[28][4]) ;
            end
            begin
              @(final_operation[28][5]) ;
            end
            begin
              @(final_operation[28][6]) ;
            end
            begin
              @(final_operation[28][7]) ;
            end
            begin
              @(final_operation[28][8]) ;
            end
            begin
              @(final_operation[28][9]) ;
            end
            begin
              @(final_operation[28][10]) ;
            end
            begin
              @(final_operation[28][11]) ;
            end
            begin
              @(final_operation[28][12]) ;
            end
            begin
              @(final_operation[28][13]) ;
            end
            begin
              @(final_operation[28][14]) ;
            end
            begin
              @(final_operation[28][15]) ;
            end
            begin
              @(final_operation[28][16]) ;
            end
            begin
              @(final_operation[28][17]) ;
            end
            begin
              @(final_operation[28][18]) ;
            end
            begin
              @(final_operation[28][19]) ;
            end
            begin
              @(final_operation[28][20]) ;
            end
            begin
              @(final_operation[28][21]) ;
            end
            begin
              @(final_operation[28][22]) ;
            end
            begin
              @(final_operation[28][23]) ;
            end
            begin
              @(final_operation[28][24]) ;
            end
            begin
              @(final_operation[28][25]) ;
            end
            begin
              @(final_operation[28][26]) ;
            end
            begin
              @(final_operation[28][27]) ;
            end
            begin
              @(final_operation[28][28]) ;
            end
            begin
              @(final_operation[28][29]) ;
            end
            begin
              @(final_operation[28][30]) ;
            end
            begin
              @(final_operation[28][31]) ;
            end

            begin
              @(final_operation[29][0]) ;
            end
            begin
              @(final_operation[29][1]) ;
            end
            begin
              @(final_operation[29][2]) ;
            end
            begin
              @(final_operation[29][3]) ;
            end
            begin
              @(final_operation[29][4]) ;
            end
            begin
              @(final_operation[29][5]) ;
            end
            begin
              @(final_operation[29][6]) ;
            end
            begin
              @(final_operation[29][7]) ;
            end
            begin
              @(final_operation[29][8]) ;
            end
            begin
              @(final_operation[29][9]) ;
            end
            begin
              @(final_operation[29][10]) ;
            end
            begin
              @(final_operation[29][11]) ;
            end
            begin
              @(final_operation[29][12]) ;
            end
            begin
              @(final_operation[29][13]) ;
            end
            begin
              @(final_operation[29][14]) ;
            end
            begin
              @(final_operation[29][15]) ;
            end
            begin
              @(final_operation[29][16]) ;
            end
            begin
              @(final_operation[29][17]) ;
            end
            begin
              @(final_operation[29][18]) ;
            end
            begin
              @(final_operation[29][19]) ;
            end
            begin
              @(final_operation[29][20]) ;
            end
            begin
              @(final_operation[29][21]) ;
            end
            begin
              @(final_operation[29][22]) ;
            end
            begin
              @(final_operation[29][23]) ;
            end
            begin
              @(final_operation[29][24]) ;
            end
            begin
              @(final_operation[29][25]) ;
            end
            begin
              @(final_operation[29][26]) ;
            end
            begin
              @(final_operation[29][27]) ;
            end
            begin
              @(final_operation[29][28]) ;
            end
            begin
              @(final_operation[29][29]) ;
            end
            begin
              @(final_operation[29][30]) ;
            end
            begin
              @(final_operation[29][31]) ;
            end

            begin
              @(final_operation[30][0]) ;
            end
            begin
              @(final_operation[30][1]) ;
            end
            begin
              @(final_operation[30][2]) ;
            end
            begin
              @(final_operation[30][3]) ;
            end
            begin
              @(final_operation[30][4]) ;
            end
            begin
              @(final_operation[30][5]) ;
            end
            begin
              @(final_operation[30][6]) ;
            end
            begin
              @(final_operation[30][7]) ;
            end
            begin
              @(final_operation[30][8]) ;
            end
            begin
              @(final_operation[30][9]) ;
            end
            begin
              @(final_operation[30][10]) ;
            end
            begin
              @(final_operation[30][11]) ;
            end
            begin
              @(final_operation[30][12]) ;
            end
            begin
              @(final_operation[30][13]) ;
            end
            begin
              @(final_operation[30][14]) ;
            end
            begin
              @(final_operation[30][15]) ;
            end
            begin
              @(final_operation[30][16]) ;
            end
            begin
              @(final_operation[30][17]) ;
            end
            begin
              @(final_operation[30][18]) ;
            end
            begin
              @(final_operation[30][19]) ;
            end
            begin
              @(final_operation[30][20]) ;
            end
            begin
              @(final_operation[30][21]) ;
            end
            begin
              @(final_operation[30][22]) ;
            end
            begin
              @(final_operation[30][23]) ;
            end
            begin
              @(final_operation[30][24]) ;
            end
            begin
              @(final_operation[30][25]) ;
            end
            begin
              @(final_operation[30][26]) ;
            end
            begin
              @(final_operation[30][27]) ;
            end
            begin
              @(final_operation[30][28]) ;
            end
            begin
              @(final_operation[30][29]) ;
            end
            begin
              @(final_operation[30][30]) ;
            end
            begin
              @(final_operation[30][31]) ;
            end

            begin
              @(final_operation[31][0]) ;
            end
            begin
              @(final_operation[31][1]) ;
            end
            begin
              @(final_operation[31][2]) ;
            end
            begin
              @(final_operation[31][3]) ;
            end
            begin
              @(final_operation[31][4]) ;
            end
            begin
              @(final_operation[31][5]) ;
            end
            begin
              @(final_operation[31][6]) ;
            end
            begin
              @(final_operation[31][7]) ;
            end
            begin
              @(final_operation[31][8]) ;
            end
            begin
              @(final_operation[31][9]) ;
            end
            begin
              @(final_operation[31][10]) ;
            end
            begin
              @(final_operation[31][11]) ;
            end
            begin
              @(final_operation[31][12]) ;
            end
            begin
              @(final_operation[31][13]) ;
            end
            begin
              @(final_operation[31][14]) ;
            end
            begin
              @(final_operation[31][15]) ;
            end
            begin
              @(final_operation[31][16]) ;
            end
            begin
              @(final_operation[31][17]) ;
            end
            begin
              @(final_operation[31][18]) ;
            end
            begin
              @(final_operation[31][19]) ;
            end
            begin
              @(final_operation[31][20]) ;
            end
            begin
              @(final_operation[31][21]) ;
            end
            begin
              @(final_operation[31][22]) ;
            end
            begin
              @(final_operation[31][23]) ;
            end
            begin
              @(final_operation[31][24]) ;
            end
            begin
              @(final_operation[31][25]) ;
            end
            begin
              @(final_operation[31][26]) ;
            end
            begin
              @(final_operation[31][27]) ;
            end
            begin
              @(final_operation[31][28]) ;
            end
            begin
              @(final_operation[31][29]) ;
            end
            begin
              @(final_operation[31][30]) ;
            end
            begin
              @(final_operation[31][31]) ;
            end

            begin
              @(final_operation[32][0]) ;
            end
            begin
              @(final_operation[32][1]) ;
            end
            begin
              @(final_operation[32][2]) ;
            end
            begin
              @(final_operation[32][3]) ;
            end
            begin
              @(final_operation[32][4]) ;
            end
            begin
              @(final_operation[32][5]) ;
            end
            begin
              @(final_operation[32][6]) ;
            end
            begin
              @(final_operation[32][7]) ;
            end
            begin
              @(final_operation[32][8]) ;
            end
            begin
              @(final_operation[32][9]) ;
            end
            begin
              @(final_operation[32][10]) ;
            end
            begin
              @(final_operation[32][11]) ;
            end
            begin
              @(final_operation[32][12]) ;
            end
            begin
              @(final_operation[32][13]) ;
            end
            begin
              @(final_operation[32][14]) ;
            end
            begin
              @(final_operation[32][15]) ;
            end
            begin
              @(final_operation[32][16]) ;
            end
            begin
              @(final_operation[32][17]) ;
            end
            begin
              @(final_operation[32][18]) ;
            end
            begin
              @(final_operation[32][19]) ;
            end
            begin
              @(final_operation[32][20]) ;
            end
            begin
              @(final_operation[32][21]) ;
            end
            begin
              @(final_operation[32][22]) ;
            end
            begin
              @(final_operation[32][23]) ;
            end
            begin
              @(final_operation[32][24]) ;
            end
            begin
              @(final_operation[32][25]) ;
            end
            begin
              @(final_operation[32][26]) ;
            end
            begin
              @(final_operation[32][27]) ;
            end
            begin
              @(final_operation[32][28]) ;
            end
            begin
              @(final_operation[32][29]) ;
            end
            begin
              @(final_operation[32][30]) ;
            end
            begin
              @(final_operation[32][31]) ;
            end

            begin
              @(final_operation[33][0]) ;
            end
            begin
              @(final_operation[33][1]) ;
            end
            begin
              @(final_operation[33][2]) ;
            end
            begin
              @(final_operation[33][3]) ;
            end
            begin
              @(final_operation[33][4]) ;
            end
            begin
              @(final_operation[33][5]) ;
            end
            begin
              @(final_operation[33][6]) ;
            end
            begin
              @(final_operation[33][7]) ;
            end
            begin
              @(final_operation[33][8]) ;
            end
            begin
              @(final_operation[33][9]) ;
            end
            begin
              @(final_operation[33][10]) ;
            end
            begin
              @(final_operation[33][11]) ;
            end
            begin
              @(final_operation[33][12]) ;
            end
            begin
              @(final_operation[33][13]) ;
            end
            begin
              @(final_operation[33][14]) ;
            end
            begin
              @(final_operation[33][15]) ;
            end
            begin
              @(final_operation[33][16]) ;
            end
            begin
              @(final_operation[33][17]) ;
            end
            begin
              @(final_operation[33][18]) ;
            end
            begin
              @(final_operation[33][19]) ;
            end
            begin
              @(final_operation[33][20]) ;
            end
            begin
              @(final_operation[33][21]) ;
            end
            begin
              @(final_operation[33][22]) ;
            end
            begin
              @(final_operation[33][23]) ;
            end
            begin
              @(final_operation[33][24]) ;
            end
            begin
              @(final_operation[33][25]) ;
            end
            begin
              @(final_operation[33][26]) ;
            end
            begin
              @(final_operation[33][27]) ;
            end
            begin
              @(final_operation[33][28]) ;
            end
            begin
              @(final_operation[33][29]) ;
            end
            begin
              @(final_operation[33][30]) ;
            end
            begin
              @(final_operation[33][31]) ;
            end

            begin
              @(final_operation[34][0]) ;
            end
            begin
              @(final_operation[34][1]) ;
            end
            begin
              @(final_operation[34][2]) ;
            end
            begin
              @(final_operation[34][3]) ;
            end
            begin
              @(final_operation[34][4]) ;
            end
            begin
              @(final_operation[34][5]) ;
            end
            begin
              @(final_operation[34][6]) ;
            end
            begin
              @(final_operation[34][7]) ;
            end
            begin
              @(final_operation[34][8]) ;
            end
            begin
              @(final_operation[34][9]) ;
            end
            begin
              @(final_operation[34][10]) ;
            end
            begin
              @(final_operation[34][11]) ;
            end
            begin
              @(final_operation[34][12]) ;
            end
            begin
              @(final_operation[34][13]) ;
            end
            begin
              @(final_operation[34][14]) ;
            end
            begin
              @(final_operation[34][15]) ;
            end
            begin
              @(final_operation[34][16]) ;
            end
            begin
              @(final_operation[34][17]) ;
            end
            begin
              @(final_operation[34][18]) ;
            end
            begin
              @(final_operation[34][19]) ;
            end
            begin
              @(final_operation[34][20]) ;
            end
            begin
              @(final_operation[34][21]) ;
            end
            begin
              @(final_operation[34][22]) ;
            end
            begin
              @(final_operation[34][23]) ;
            end
            begin
              @(final_operation[34][24]) ;
            end
            begin
              @(final_operation[34][25]) ;
            end
            begin
              @(final_operation[34][26]) ;
            end
            begin
              @(final_operation[34][27]) ;
            end
            begin
              @(final_operation[34][28]) ;
            end
            begin
              @(final_operation[34][29]) ;
            end
            begin
              @(final_operation[34][30]) ;
            end
            begin
              @(final_operation[34][31]) ;
            end

            begin
              @(final_operation[35][0]) ;
            end
            begin
              @(final_operation[35][1]) ;
            end
            begin
              @(final_operation[35][2]) ;
            end
            begin
              @(final_operation[35][3]) ;
            end
            begin
              @(final_operation[35][4]) ;
            end
            begin
              @(final_operation[35][5]) ;
            end
            begin
              @(final_operation[35][6]) ;
            end
            begin
              @(final_operation[35][7]) ;
            end
            begin
              @(final_operation[35][8]) ;
            end
            begin
              @(final_operation[35][9]) ;
            end
            begin
              @(final_operation[35][10]) ;
            end
            begin
              @(final_operation[35][11]) ;
            end
            begin
              @(final_operation[35][12]) ;
            end
            begin
              @(final_operation[35][13]) ;
            end
            begin
              @(final_operation[35][14]) ;
            end
            begin
              @(final_operation[35][15]) ;
            end
            begin
              @(final_operation[35][16]) ;
            end
            begin
              @(final_operation[35][17]) ;
            end
            begin
              @(final_operation[35][18]) ;
            end
            begin
              @(final_operation[35][19]) ;
            end
            begin
              @(final_operation[35][20]) ;
            end
            begin
              @(final_operation[35][21]) ;
            end
            begin
              @(final_operation[35][22]) ;
            end
            begin
              @(final_operation[35][23]) ;
            end
            begin
              @(final_operation[35][24]) ;
            end
            begin
              @(final_operation[35][25]) ;
            end
            begin
              @(final_operation[35][26]) ;
            end
            begin
              @(final_operation[35][27]) ;
            end
            begin
              @(final_operation[35][28]) ;
            end
            begin
              @(final_operation[35][29]) ;
            end
            begin
              @(final_operation[35][30]) ;
            end
            begin
              @(final_operation[35][31]) ;
            end

            begin
              @(final_operation[36][0]) ;
            end
            begin
              @(final_operation[36][1]) ;
            end
            begin
              @(final_operation[36][2]) ;
            end
            begin
              @(final_operation[36][3]) ;
            end
            begin
              @(final_operation[36][4]) ;
            end
            begin
              @(final_operation[36][5]) ;
            end
            begin
              @(final_operation[36][6]) ;
            end
            begin
              @(final_operation[36][7]) ;
            end
            begin
              @(final_operation[36][8]) ;
            end
            begin
              @(final_operation[36][9]) ;
            end
            begin
              @(final_operation[36][10]) ;
            end
            begin
              @(final_operation[36][11]) ;
            end
            begin
              @(final_operation[36][12]) ;
            end
            begin
              @(final_operation[36][13]) ;
            end
            begin
              @(final_operation[36][14]) ;
            end
            begin
              @(final_operation[36][15]) ;
            end
            begin
              @(final_operation[36][16]) ;
            end
            begin
              @(final_operation[36][17]) ;
            end
            begin
              @(final_operation[36][18]) ;
            end
            begin
              @(final_operation[36][19]) ;
            end
            begin
              @(final_operation[36][20]) ;
            end
            begin
              @(final_operation[36][21]) ;
            end
            begin
              @(final_operation[36][22]) ;
            end
            begin
              @(final_operation[36][23]) ;
            end
            begin
              @(final_operation[36][24]) ;
            end
            begin
              @(final_operation[36][25]) ;
            end
            begin
              @(final_operation[36][26]) ;
            end
            begin
              @(final_operation[36][27]) ;
            end
            begin
              @(final_operation[36][28]) ;
            end
            begin
              @(final_operation[36][29]) ;
            end
            begin
              @(final_operation[36][30]) ;
            end
            begin
              @(final_operation[36][31]) ;
            end

            begin
              @(final_operation[37][0]) ;
            end
            begin
              @(final_operation[37][1]) ;
            end
            begin
              @(final_operation[37][2]) ;
            end
            begin
              @(final_operation[37][3]) ;
            end
            begin
              @(final_operation[37][4]) ;
            end
            begin
              @(final_operation[37][5]) ;
            end
            begin
              @(final_operation[37][6]) ;
            end
            begin
              @(final_operation[37][7]) ;
            end
            begin
              @(final_operation[37][8]) ;
            end
            begin
              @(final_operation[37][9]) ;
            end
            begin
              @(final_operation[37][10]) ;
            end
            begin
              @(final_operation[37][11]) ;
            end
            begin
              @(final_operation[37][12]) ;
            end
            begin
              @(final_operation[37][13]) ;
            end
            begin
              @(final_operation[37][14]) ;
            end
            begin
              @(final_operation[37][15]) ;
            end
            begin
              @(final_operation[37][16]) ;
            end
            begin
              @(final_operation[37][17]) ;
            end
            begin
              @(final_operation[37][18]) ;
            end
            begin
              @(final_operation[37][19]) ;
            end
            begin
              @(final_operation[37][20]) ;
            end
            begin
              @(final_operation[37][21]) ;
            end
            begin
              @(final_operation[37][22]) ;
            end
            begin
              @(final_operation[37][23]) ;
            end
            begin
              @(final_operation[37][24]) ;
            end
            begin
              @(final_operation[37][25]) ;
            end
            begin
              @(final_operation[37][26]) ;
            end
            begin
              @(final_operation[37][27]) ;
            end
            begin
              @(final_operation[37][28]) ;
            end
            begin
              @(final_operation[37][29]) ;
            end
            begin
              @(final_operation[37][30]) ;
            end
            begin
              @(final_operation[37][31]) ;
            end

            begin
              @(final_operation[38][0]) ;
            end
            begin
              @(final_operation[38][1]) ;
            end
            begin
              @(final_operation[38][2]) ;
            end
            begin
              @(final_operation[38][3]) ;
            end
            begin
              @(final_operation[38][4]) ;
            end
            begin
              @(final_operation[38][5]) ;
            end
            begin
              @(final_operation[38][6]) ;
            end
            begin
              @(final_operation[38][7]) ;
            end
            begin
              @(final_operation[38][8]) ;
            end
            begin
              @(final_operation[38][9]) ;
            end
            begin
              @(final_operation[38][10]) ;
            end
            begin
              @(final_operation[38][11]) ;
            end
            begin
              @(final_operation[38][12]) ;
            end
            begin
              @(final_operation[38][13]) ;
            end
            begin
              @(final_operation[38][14]) ;
            end
            begin
              @(final_operation[38][15]) ;
            end
            begin
              @(final_operation[38][16]) ;
            end
            begin
              @(final_operation[38][17]) ;
            end
            begin
              @(final_operation[38][18]) ;
            end
            begin
              @(final_operation[38][19]) ;
            end
            begin
              @(final_operation[38][20]) ;
            end
            begin
              @(final_operation[38][21]) ;
            end
            begin
              @(final_operation[38][22]) ;
            end
            begin
              @(final_operation[38][23]) ;
            end
            begin
              @(final_operation[38][24]) ;
            end
            begin
              @(final_operation[38][25]) ;
            end
            begin
              @(final_operation[38][26]) ;
            end
            begin
              @(final_operation[38][27]) ;
            end
            begin
              @(final_operation[38][28]) ;
            end
            begin
              @(final_operation[38][29]) ;
            end
            begin
              @(final_operation[38][30]) ;
            end
            begin
              @(final_operation[38][31]) ;
            end

            begin
              @(final_operation[39][0]) ;
            end
            begin
              @(final_operation[39][1]) ;
            end
            begin
              @(final_operation[39][2]) ;
            end
            begin
              @(final_operation[39][3]) ;
            end
            begin
              @(final_operation[39][4]) ;
            end
            begin
              @(final_operation[39][5]) ;
            end
            begin
              @(final_operation[39][6]) ;
            end
            begin
              @(final_operation[39][7]) ;
            end
            begin
              @(final_operation[39][8]) ;
            end
            begin
              @(final_operation[39][9]) ;
            end
            begin
              @(final_operation[39][10]) ;
            end
            begin
              @(final_operation[39][11]) ;
            end
            begin
              @(final_operation[39][12]) ;
            end
            begin
              @(final_operation[39][13]) ;
            end
            begin
              @(final_operation[39][14]) ;
            end
            begin
              @(final_operation[39][15]) ;
            end
            begin
              @(final_operation[39][16]) ;
            end
            begin
              @(final_operation[39][17]) ;
            end
            begin
              @(final_operation[39][18]) ;
            end
            begin
              @(final_operation[39][19]) ;
            end
            begin
              @(final_operation[39][20]) ;
            end
            begin
              @(final_operation[39][21]) ;
            end
            begin
              @(final_operation[39][22]) ;
            end
            begin
              @(final_operation[39][23]) ;
            end
            begin
              @(final_operation[39][24]) ;
            end
            begin
              @(final_operation[39][25]) ;
            end
            begin
              @(final_operation[39][26]) ;
            end
            begin
              @(final_operation[39][27]) ;
            end
            begin
              @(final_operation[39][28]) ;
            end
            begin
              @(final_operation[39][29]) ;
            end
            begin
              @(final_operation[39][30]) ;
            end
            begin
              @(final_operation[39][31]) ;
            end

            begin
              @(final_operation[40][0]) ;
            end
            begin
              @(final_operation[40][1]) ;
            end
            begin
              @(final_operation[40][2]) ;
            end
            begin
              @(final_operation[40][3]) ;
            end
            begin
              @(final_operation[40][4]) ;
            end
            begin
              @(final_operation[40][5]) ;
            end
            begin
              @(final_operation[40][6]) ;
            end
            begin
              @(final_operation[40][7]) ;
            end
            begin
              @(final_operation[40][8]) ;
            end
            begin
              @(final_operation[40][9]) ;
            end
            begin
              @(final_operation[40][10]) ;
            end
            begin
              @(final_operation[40][11]) ;
            end
            begin
              @(final_operation[40][12]) ;
            end
            begin
              @(final_operation[40][13]) ;
            end
            begin
              @(final_operation[40][14]) ;
            end
            begin
              @(final_operation[40][15]) ;
            end
            begin
              @(final_operation[40][16]) ;
            end
            begin
              @(final_operation[40][17]) ;
            end
            begin
              @(final_operation[40][18]) ;
            end
            begin
              @(final_operation[40][19]) ;
            end
            begin
              @(final_operation[40][20]) ;
            end
            begin
              @(final_operation[40][21]) ;
            end
            begin
              @(final_operation[40][22]) ;
            end
            begin
              @(final_operation[40][23]) ;
            end
            begin
              @(final_operation[40][24]) ;
            end
            begin
              @(final_operation[40][25]) ;
            end
            begin
              @(final_operation[40][26]) ;
            end
            begin
              @(final_operation[40][27]) ;
            end
            begin
              @(final_operation[40][28]) ;
            end
            begin
              @(final_operation[40][29]) ;
            end
            begin
              @(final_operation[40][30]) ;
            end
            begin
              @(final_operation[40][31]) ;
            end

            begin
              @(final_operation[41][0]) ;
            end
            begin
              @(final_operation[41][1]) ;
            end
            begin
              @(final_operation[41][2]) ;
            end
            begin
              @(final_operation[41][3]) ;
            end
            begin
              @(final_operation[41][4]) ;
            end
            begin
              @(final_operation[41][5]) ;
            end
            begin
              @(final_operation[41][6]) ;
            end
            begin
              @(final_operation[41][7]) ;
            end
            begin
              @(final_operation[41][8]) ;
            end
            begin
              @(final_operation[41][9]) ;
            end
            begin
              @(final_operation[41][10]) ;
            end
            begin
              @(final_operation[41][11]) ;
            end
            begin
              @(final_operation[41][12]) ;
            end
            begin
              @(final_operation[41][13]) ;
            end
            begin
              @(final_operation[41][14]) ;
            end
            begin
              @(final_operation[41][15]) ;
            end
            begin
              @(final_operation[41][16]) ;
            end
            begin
              @(final_operation[41][17]) ;
            end
            begin
              @(final_operation[41][18]) ;
            end
            begin
              @(final_operation[41][19]) ;
            end
            begin
              @(final_operation[41][20]) ;
            end
            begin
              @(final_operation[41][21]) ;
            end
            begin
              @(final_operation[41][22]) ;
            end
            begin
              @(final_operation[41][23]) ;
            end
            begin
              @(final_operation[41][24]) ;
            end
            begin
              @(final_operation[41][25]) ;
            end
            begin
              @(final_operation[41][26]) ;
            end
            begin
              @(final_operation[41][27]) ;
            end
            begin
              @(final_operation[41][28]) ;
            end
            begin
              @(final_operation[41][29]) ;
            end
            begin
              @(final_operation[41][30]) ;
            end
            begin
              @(final_operation[41][31]) ;
            end

            begin
              @(final_operation[42][0]) ;
            end
            begin
              @(final_operation[42][1]) ;
            end
            begin
              @(final_operation[42][2]) ;
            end
            begin
              @(final_operation[42][3]) ;
            end
            begin
              @(final_operation[42][4]) ;
            end
            begin
              @(final_operation[42][5]) ;
            end
            begin
              @(final_operation[42][6]) ;
            end
            begin
              @(final_operation[42][7]) ;
            end
            begin
              @(final_operation[42][8]) ;
            end
            begin
              @(final_operation[42][9]) ;
            end
            begin
              @(final_operation[42][10]) ;
            end
            begin
              @(final_operation[42][11]) ;
            end
            begin
              @(final_operation[42][12]) ;
            end
            begin
              @(final_operation[42][13]) ;
            end
            begin
              @(final_operation[42][14]) ;
            end
            begin
              @(final_operation[42][15]) ;
            end
            begin
              @(final_operation[42][16]) ;
            end
            begin
              @(final_operation[42][17]) ;
            end
            begin
              @(final_operation[42][18]) ;
            end
            begin
              @(final_operation[42][19]) ;
            end
            begin
              @(final_operation[42][20]) ;
            end
            begin
              @(final_operation[42][21]) ;
            end
            begin
              @(final_operation[42][22]) ;
            end
            begin
              @(final_operation[42][23]) ;
            end
            begin
              @(final_operation[42][24]) ;
            end
            begin
              @(final_operation[42][25]) ;
            end
            begin
              @(final_operation[42][26]) ;
            end
            begin
              @(final_operation[42][27]) ;
            end
            begin
              @(final_operation[42][28]) ;
            end
            begin
              @(final_operation[42][29]) ;
            end
            begin
              @(final_operation[42][30]) ;
            end
            begin
              @(final_operation[42][31]) ;
            end

            begin
              @(final_operation[43][0]) ;
            end
            begin
              @(final_operation[43][1]) ;
            end
            begin
              @(final_operation[43][2]) ;
            end
            begin
              @(final_operation[43][3]) ;
            end
            begin
              @(final_operation[43][4]) ;
            end
            begin
              @(final_operation[43][5]) ;
            end
            begin
              @(final_operation[43][6]) ;
            end
            begin
              @(final_operation[43][7]) ;
            end
            begin
              @(final_operation[43][8]) ;
            end
            begin
              @(final_operation[43][9]) ;
            end
            begin
              @(final_operation[43][10]) ;
            end
            begin
              @(final_operation[43][11]) ;
            end
            begin
              @(final_operation[43][12]) ;
            end
            begin
              @(final_operation[43][13]) ;
            end
            begin
              @(final_operation[43][14]) ;
            end
            begin
              @(final_operation[43][15]) ;
            end
            begin
              @(final_operation[43][16]) ;
            end
            begin
              @(final_operation[43][17]) ;
            end
            begin
              @(final_operation[43][18]) ;
            end
            begin
              @(final_operation[43][19]) ;
            end
            begin
              @(final_operation[43][20]) ;
            end
            begin
              @(final_operation[43][21]) ;
            end
            begin
              @(final_operation[43][22]) ;
            end
            begin
              @(final_operation[43][23]) ;
            end
            begin
              @(final_operation[43][24]) ;
            end
            begin
              @(final_operation[43][25]) ;
            end
            begin
              @(final_operation[43][26]) ;
            end
            begin
              @(final_operation[43][27]) ;
            end
            begin
              @(final_operation[43][28]) ;
            end
            begin
              @(final_operation[43][29]) ;
            end
            begin
              @(final_operation[43][30]) ;
            end
            begin
              @(final_operation[43][31]) ;
            end

            begin
              @(final_operation[44][0]) ;
            end
            begin
              @(final_operation[44][1]) ;
            end
            begin
              @(final_operation[44][2]) ;
            end
            begin
              @(final_operation[44][3]) ;
            end
            begin
              @(final_operation[44][4]) ;
            end
            begin
              @(final_operation[44][5]) ;
            end
            begin
              @(final_operation[44][6]) ;
            end
            begin
              @(final_operation[44][7]) ;
            end
            begin
              @(final_operation[44][8]) ;
            end
            begin
              @(final_operation[44][9]) ;
            end
            begin
              @(final_operation[44][10]) ;
            end
            begin
              @(final_operation[44][11]) ;
            end
            begin
              @(final_operation[44][12]) ;
            end
            begin
              @(final_operation[44][13]) ;
            end
            begin
              @(final_operation[44][14]) ;
            end
            begin
              @(final_operation[44][15]) ;
            end
            begin
              @(final_operation[44][16]) ;
            end
            begin
              @(final_operation[44][17]) ;
            end
            begin
              @(final_operation[44][18]) ;
            end
            begin
              @(final_operation[44][19]) ;
            end
            begin
              @(final_operation[44][20]) ;
            end
            begin
              @(final_operation[44][21]) ;
            end
            begin
              @(final_operation[44][22]) ;
            end
            begin
              @(final_operation[44][23]) ;
            end
            begin
              @(final_operation[44][24]) ;
            end
            begin
              @(final_operation[44][25]) ;
            end
            begin
              @(final_operation[44][26]) ;
            end
            begin
              @(final_operation[44][27]) ;
            end
            begin
              @(final_operation[44][28]) ;
            end
            begin
              @(final_operation[44][29]) ;
            end
            begin
              @(final_operation[44][30]) ;
            end
            begin
              @(final_operation[44][31]) ;
            end

            begin
              @(final_operation[45][0]) ;
            end
            begin
              @(final_operation[45][1]) ;
            end
            begin
              @(final_operation[45][2]) ;
            end
            begin
              @(final_operation[45][3]) ;
            end
            begin
              @(final_operation[45][4]) ;
            end
            begin
              @(final_operation[45][5]) ;
            end
            begin
              @(final_operation[45][6]) ;
            end
            begin
              @(final_operation[45][7]) ;
            end
            begin
              @(final_operation[45][8]) ;
            end
            begin
              @(final_operation[45][9]) ;
            end
            begin
              @(final_operation[45][10]) ;
            end
            begin
              @(final_operation[45][11]) ;
            end
            begin
              @(final_operation[45][12]) ;
            end
            begin
              @(final_operation[45][13]) ;
            end
            begin
              @(final_operation[45][14]) ;
            end
            begin
              @(final_operation[45][15]) ;
            end
            begin
              @(final_operation[45][16]) ;
            end
            begin
              @(final_operation[45][17]) ;
            end
            begin
              @(final_operation[45][18]) ;
            end
            begin
              @(final_operation[45][19]) ;
            end
            begin
              @(final_operation[45][20]) ;
            end
            begin
              @(final_operation[45][21]) ;
            end
            begin
              @(final_operation[45][22]) ;
            end
            begin
              @(final_operation[45][23]) ;
            end
            begin
              @(final_operation[45][24]) ;
            end
            begin
              @(final_operation[45][25]) ;
            end
            begin
              @(final_operation[45][26]) ;
            end
            begin
              @(final_operation[45][27]) ;
            end
            begin
              @(final_operation[45][28]) ;
            end
            begin
              @(final_operation[45][29]) ;
            end
            begin
              @(final_operation[45][30]) ;
            end
            begin
              @(final_operation[45][31]) ;
            end

            begin
              @(final_operation[46][0]) ;
            end
            begin
              @(final_operation[46][1]) ;
            end
            begin
              @(final_operation[46][2]) ;
            end
            begin
              @(final_operation[46][3]) ;
            end
            begin
              @(final_operation[46][4]) ;
            end
            begin
              @(final_operation[46][5]) ;
            end
            begin
              @(final_operation[46][6]) ;
            end
            begin
              @(final_operation[46][7]) ;
            end
            begin
              @(final_operation[46][8]) ;
            end
            begin
              @(final_operation[46][9]) ;
            end
            begin
              @(final_operation[46][10]) ;
            end
            begin
              @(final_operation[46][11]) ;
            end
            begin
              @(final_operation[46][12]) ;
            end
            begin
              @(final_operation[46][13]) ;
            end
            begin
              @(final_operation[46][14]) ;
            end
            begin
              @(final_operation[46][15]) ;
            end
            begin
              @(final_operation[46][16]) ;
            end
            begin
              @(final_operation[46][17]) ;
            end
            begin
              @(final_operation[46][18]) ;
            end
            begin
              @(final_operation[46][19]) ;
            end
            begin
              @(final_operation[46][20]) ;
            end
            begin
              @(final_operation[46][21]) ;
            end
            begin
              @(final_operation[46][22]) ;
            end
            begin
              @(final_operation[46][23]) ;
            end
            begin
              @(final_operation[46][24]) ;
            end
            begin
              @(final_operation[46][25]) ;
            end
            begin
              @(final_operation[46][26]) ;
            end
            begin
              @(final_operation[46][27]) ;
            end
            begin
              @(final_operation[46][28]) ;
            end
            begin
              @(final_operation[46][29]) ;
            end
            begin
              @(final_operation[46][30]) ;
            end
            begin
              @(final_operation[46][31]) ;
            end

            begin
              @(final_operation[47][0]) ;
            end
            begin
              @(final_operation[47][1]) ;
            end
            begin
              @(final_operation[47][2]) ;
            end
            begin
              @(final_operation[47][3]) ;
            end
            begin
              @(final_operation[47][4]) ;
            end
            begin
              @(final_operation[47][5]) ;
            end
            begin
              @(final_operation[47][6]) ;
            end
            begin
              @(final_operation[47][7]) ;
            end
            begin
              @(final_operation[47][8]) ;
            end
            begin
              @(final_operation[47][9]) ;
            end
            begin
              @(final_operation[47][10]) ;
            end
            begin
              @(final_operation[47][11]) ;
            end
            begin
              @(final_operation[47][12]) ;
            end
            begin
              @(final_operation[47][13]) ;
            end
            begin
              @(final_operation[47][14]) ;
            end
            begin
              @(final_operation[47][15]) ;
            end
            begin
              @(final_operation[47][16]) ;
            end
            begin
              @(final_operation[47][17]) ;
            end
            begin
              @(final_operation[47][18]) ;
            end
            begin
              @(final_operation[47][19]) ;
            end
            begin
              @(final_operation[47][20]) ;
            end
            begin
              @(final_operation[47][21]) ;
            end
            begin
              @(final_operation[47][22]) ;
            end
            begin
              @(final_operation[47][23]) ;
            end
            begin
              @(final_operation[47][24]) ;
            end
            begin
              @(final_operation[47][25]) ;
            end
            begin
              @(final_operation[47][26]) ;
            end
            begin
              @(final_operation[47][27]) ;
            end
            begin
              @(final_operation[47][28]) ;
            end
            begin
              @(final_operation[47][29]) ;
            end
            begin
              @(final_operation[47][30]) ;
            end
            begin
              @(final_operation[47][31]) ;
            end

            begin
              @(final_operation[48][0]) ;
            end
            begin
              @(final_operation[48][1]) ;
            end
            begin
              @(final_operation[48][2]) ;
            end
            begin
              @(final_operation[48][3]) ;
            end
            begin
              @(final_operation[48][4]) ;
            end
            begin
              @(final_operation[48][5]) ;
            end
            begin
              @(final_operation[48][6]) ;
            end
            begin
              @(final_operation[48][7]) ;
            end
            begin
              @(final_operation[48][8]) ;
            end
            begin
              @(final_operation[48][9]) ;
            end
            begin
              @(final_operation[48][10]) ;
            end
            begin
              @(final_operation[48][11]) ;
            end
            begin
              @(final_operation[48][12]) ;
            end
            begin
              @(final_operation[48][13]) ;
            end
            begin
              @(final_operation[48][14]) ;
            end
            begin
              @(final_operation[48][15]) ;
            end
            begin
              @(final_operation[48][16]) ;
            end
            begin
              @(final_operation[48][17]) ;
            end
            begin
              @(final_operation[48][18]) ;
            end
            begin
              @(final_operation[48][19]) ;
            end
            begin
              @(final_operation[48][20]) ;
            end
            begin
              @(final_operation[48][21]) ;
            end
            begin
              @(final_operation[48][22]) ;
            end
            begin
              @(final_operation[48][23]) ;
            end
            begin
              @(final_operation[48][24]) ;
            end
            begin
              @(final_operation[48][25]) ;
            end
            begin
              @(final_operation[48][26]) ;
            end
            begin
              @(final_operation[48][27]) ;
            end
            begin
              @(final_operation[48][28]) ;
            end
            begin
              @(final_operation[48][29]) ;
            end
            begin
              @(final_operation[48][30]) ;
            end
            begin
              @(final_operation[48][31]) ;
            end

            begin
              @(final_operation[49][0]) ;
            end
            begin
              @(final_operation[49][1]) ;
            end
            begin
              @(final_operation[49][2]) ;
            end
            begin
              @(final_operation[49][3]) ;
            end
            begin
              @(final_operation[49][4]) ;
            end
            begin
              @(final_operation[49][5]) ;
            end
            begin
              @(final_operation[49][6]) ;
            end
            begin
              @(final_operation[49][7]) ;
            end
            begin
              @(final_operation[49][8]) ;
            end
            begin
              @(final_operation[49][9]) ;
            end
            begin
              @(final_operation[49][10]) ;
            end
            begin
              @(final_operation[49][11]) ;
            end
            begin
              @(final_operation[49][12]) ;
            end
            begin
              @(final_operation[49][13]) ;
            end
            begin
              @(final_operation[49][14]) ;
            end
            begin
              @(final_operation[49][15]) ;
            end
            begin
              @(final_operation[49][16]) ;
            end
            begin
              @(final_operation[49][17]) ;
            end
            begin
              @(final_operation[49][18]) ;
            end
            begin
              @(final_operation[49][19]) ;
            end
            begin
              @(final_operation[49][20]) ;
            end
            begin
              @(final_operation[49][21]) ;
            end
            begin
              @(final_operation[49][22]) ;
            end
            begin
              @(final_operation[49][23]) ;
            end
            begin
              @(final_operation[49][24]) ;
            end
            begin
              @(final_operation[49][25]) ;
            end
            begin
              @(final_operation[49][26]) ;
            end
            begin
              @(final_operation[49][27]) ;
            end
            begin
              @(final_operation[49][28]) ;
            end
            begin
              @(final_operation[49][29]) ;
            end
            begin
              @(final_operation[49][30]) ;
            end
            begin
              @(final_operation[49][31]) ;
            end

            begin
              @(final_operation[50][0]) ;
            end
            begin
              @(final_operation[50][1]) ;
            end
            begin
              @(final_operation[50][2]) ;
            end
            begin
              @(final_operation[50][3]) ;
            end
            begin
              @(final_operation[50][4]) ;
            end
            begin
              @(final_operation[50][5]) ;
            end
            begin
              @(final_operation[50][6]) ;
            end
            begin
              @(final_operation[50][7]) ;
            end
            begin
              @(final_operation[50][8]) ;
            end
            begin
              @(final_operation[50][9]) ;
            end
            begin
              @(final_operation[50][10]) ;
            end
            begin
              @(final_operation[50][11]) ;
            end
            begin
              @(final_operation[50][12]) ;
            end
            begin
              @(final_operation[50][13]) ;
            end
            begin
              @(final_operation[50][14]) ;
            end
            begin
              @(final_operation[50][15]) ;
            end
            begin
              @(final_operation[50][16]) ;
            end
            begin
              @(final_operation[50][17]) ;
            end
            begin
              @(final_operation[50][18]) ;
            end
            begin
              @(final_operation[50][19]) ;
            end
            begin
              @(final_operation[50][20]) ;
            end
            begin
              @(final_operation[50][21]) ;
            end
            begin
              @(final_operation[50][22]) ;
            end
            begin
              @(final_operation[50][23]) ;
            end
            begin
              @(final_operation[50][24]) ;
            end
            begin
              @(final_operation[50][25]) ;
            end
            begin
              @(final_operation[50][26]) ;
            end
            begin
              @(final_operation[50][27]) ;
            end
            begin
              @(final_operation[50][28]) ;
            end
            begin
              @(final_operation[50][29]) ;
            end
            begin
              @(final_operation[50][30]) ;
            end
            begin
              @(final_operation[50][31]) ;
            end

            begin
              @(final_operation[51][0]) ;
            end
            begin
              @(final_operation[51][1]) ;
            end
            begin
              @(final_operation[51][2]) ;
            end
            begin
              @(final_operation[51][3]) ;
            end
            begin
              @(final_operation[51][4]) ;
            end
            begin
              @(final_operation[51][5]) ;
            end
            begin
              @(final_operation[51][6]) ;
            end
            begin
              @(final_operation[51][7]) ;
            end
            begin
              @(final_operation[51][8]) ;
            end
            begin
              @(final_operation[51][9]) ;
            end
            begin
              @(final_operation[51][10]) ;
            end
            begin
              @(final_operation[51][11]) ;
            end
            begin
              @(final_operation[51][12]) ;
            end
            begin
              @(final_operation[51][13]) ;
            end
            begin
              @(final_operation[51][14]) ;
            end
            begin
              @(final_operation[51][15]) ;
            end
            begin
              @(final_operation[51][16]) ;
            end
            begin
              @(final_operation[51][17]) ;
            end
            begin
              @(final_operation[51][18]) ;
            end
            begin
              @(final_operation[51][19]) ;
            end
            begin
              @(final_operation[51][20]) ;
            end
            begin
              @(final_operation[51][21]) ;
            end
            begin
              @(final_operation[51][22]) ;
            end
            begin
              @(final_operation[51][23]) ;
            end
            begin
              @(final_operation[51][24]) ;
            end
            begin
              @(final_operation[51][25]) ;
            end
            begin
              @(final_operation[51][26]) ;
            end
            begin
              @(final_operation[51][27]) ;
            end
            begin
              @(final_operation[51][28]) ;
            end
            begin
              @(final_operation[51][29]) ;
            end
            begin
              @(final_operation[51][30]) ;
            end
            begin
              @(final_operation[51][31]) ;
            end

            begin
              @(final_operation[52][0]) ;
            end
            begin
              @(final_operation[52][1]) ;
            end
            begin
              @(final_operation[52][2]) ;
            end
            begin
              @(final_operation[52][3]) ;
            end
            begin
              @(final_operation[52][4]) ;
            end
            begin
              @(final_operation[52][5]) ;
            end
            begin
              @(final_operation[52][6]) ;
            end
            begin
              @(final_operation[52][7]) ;
            end
            begin
              @(final_operation[52][8]) ;
            end
            begin
              @(final_operation[52][9]) ;
            end
            begin
              @(final_operation[52][10]) ;
            end
            begin
              @(final_operation[52][11]) ;
            end
            begin
              @(final_operation[52][12]) ;
            end
            begin
              @(final_operation[52][13]) ;
            end
            begin
              @(final_operation[52][14]) ;
            end
            begin
              @(final_operation[52][15]) ;
            end
            begin
              @(final_operation[52][16]) ;
            end
            begin
              @(final_operation[52][17]) ;
            end
            begin
              @(final_operation[52][18]) ;
            end
            begin
              @(final_operation[52][19]) ;
            end
            begin
              @(final_operation[52][20]) ;
            end
            begin
              @(final_operation[52][21]) ;
            end
            begin
              @(final_operation[52][22]) ;
            end
            begin
              @(final_operation[52][23]) ;
            end
            begin
              @(final_operation[52][24]) ;
            end
            begin
              @(final_operation[52][25]) ;
            end
            begin
              @(final_operation[52][26]) ;
            end
            begin
              @(final_operation[52][27]) ;
            end
            begin
              @(final_operation[52][28]) ;
            end
            begin
              @(final_operation[52][29]) ;
            end
            begin
              @(final_operation[52][30]) ;
            end
            begin
              @(final_operation[52][31]) ;
            end

            begin
              @(final_operation[53][0]) ;
            end
            begin
              @(final_operation[53][1]) ;
            end
            begin
              @(final_operation[53][2]) ;
            end
            begin
              @(final_operation[53][3]) ;
            end
            begin
              @(final_operation[53][4]) ;
            end
            begin
              @(final_operation[53][5]) ;
            end
            begin
              @(final_operation[53][6]) ;
            end
            begin
              @(final_operation[53][7]) ;
            end
            begin
              @(final_operation[53][8]) ;
            end
            begin
              @(final_operation[53][9]) ;
            end
            begin
              @(final_operation[53][10]) ;
            end
            begin
              @(final_operation[53][11]) ;
            end
            begin
              @(final_operation[53][12]) ;
            end
            begin
              @(final_operation[53][13]) ;
            end
            begin
              @(final_operation[53][14]) ;
            end
            begin
              @(final_operation[53][15]) ;
            end
            begin
              @(final_operation[53][16]) ;
            end
            begin
              @(final_operation[53][17]) ;
            end
            begin
              @(final_operation[53][18]) ;
            end
            begin
              @(final_operation[53][19]) ;
            end
            begin
              @(final_operation[53][20]) ;
            end
            begin
              @(final_operation[53][21]) ;
            end
            begin
              @(final_operation[53][22]) ;
            end
            begin
              @(final_operation[53][23]) ;
            end
            begin
              @(final_operation[53][24]) ;
            end
            begin
              @(final_operation[53][25]) ;
            end
            begin
              @(final_operation[53][26]) ;
            end
            begin
              @(final_operation[53][27]) ;
            end
            begin
              @(final_operation[53][28]) ;
            end
            begin
              @(final_operation[53][29]) ;
            end
            begin
              @(final_operation[53][30]) ;
            end
            begin
              @(final_operation[53][31]) ;
            end

            begin
              @(final_operation[54][0]) ;
            end
            begin
              @(final_operation[54][1]) ;
            end
            begin
              @(final_operation[54][2]) ;
            end
            begin
              @(final_operation[54][3]) ;
            end
            begin
              @(final_operation[54][4]) ;
            end
            begin
              @(final_operation[54][5]) ;
            end
            begin
              @(final_operation[54][6]) ;
            end
            begin
              @(final_operation[54][7]) ;
            end
            begin
              @(final_operation[54][8]) ;
            end
            begin
              @(final_operation[54][9]) ;
            end
            begin
              @(final_operation[54][10]) ;
            end
            begin
              @(final_operation[54][11]) ;
            end
            begin
              @(final_operation[54][12]) ;
            end
            begin
              @(final_operation[54][13]) ;
            end
            begin
              @(final_operation[54][14]) ;
            end
            begin
              @(final_operation[54][15]) ;
            end
            begin
              @(final_operation[54][16]) ;
            end
            begin
              @(final_operation[54][17]) ;
            end
            begin
              @(final_operation[54][18]) ;
            end
            begin
              @(final_operation[54][19]) ;
            end
            begin
              @(final_operation[54][20]) ;
            end
            begin
              @(final_operation[54][21]) ;
            end
            begin
              @(final_operation[54][22]) ;
            end
            begin
              @(final_operation[54][23]) ;
            end
            begin
              @(final_operation[54][24]) ;
            end
            begin
              @(final_operation[54][25]) ;
            end
            begin
              @(final_operation[54][26]) ;
            end
            begin
              @(final_operation[54][27]) ;
            end
            begin
              @(final_operation[54][28]) ;
            end
            begin
              @(final_operation[54][29]) ;
            end
            begin
              @(final_operation[54][30]) ;
            end
            begin
              @(final_operation[54][31]) ;
            end

            begin
              @(final_operation[55][0]) ;
            end
            begin
              @(final_operation[55][1]) ;
            end
            begin
              @(final_operation[55][2]) ;
            end
            begin
              @(final_operation[55][3]) ;
            end
            begin
              @(final_operation[55][4]) ;
            end
            begin
              @(final_operation[55][5]) ;
            end
            begin
              @(final_operation[55][6]) ;
            end
            begin
              @(final_operation[55][7]) ;
            end
            begin
              @(final_operation[55][8]) ;
            end
            begin
              @(final_operation[55][9]) ;
            end
            begin
              @(final_operation[55][10]) ;
            end
            begin
              @(final_operation[55][11]) ;
            end
            begin
              @(final_operation[55][12]) ;
            end
            begin
              @(final_operation[55][13]) ;
            end
            begin
              @(final_operation[55][14]) ;
            end
            begin
              @(final_operation[55][15]) ;
            end
            begin
              @(final_operation[55][16]) ;
            end
            begin
              @(final_operation[55][17]) ;
            end
            begin
              @(final_operation[55][18]) ;
            end
            begin
              @(final_operation[55][19]) ;
            end
            begin
              @(final_operation[55][20]) ;
            end
            begin
              @(final_operation[55][21]) ;
            end
            begin
              @(final_operation[55][22]) ;
            end
            begin
              @(final_operation[55][23]) ;
            end
            begin
              @(final_operation[55][24]) ;
            end
            begin
              @(final_operation[55][25]) ;
            end
            begin
              @(final_operation[55][26]) ;
            end
            begin
              @(final_operation[55][27]) ;
            end
            begin
              @(final_operation[55][28]) ;
            end
            begin
              @(final_operation[55][29]) ;
            end
            begin
              @(final_operation[55][30]) ;
            end
            begin
              @(final_operation[55][31]) ;
            end

            begin
              @(final_operation[56][0]) ;
            end
            begin
              @(final_operation[56][1]) ;
            end
            begin
              @(final_operation[56][2]) ;
            end
            begin
              @(final_operation[56][3]) ;
            end
            begin
              @(final_operation[56][4]) ;
            end
            begin
              @(final_operation[56][5]) ;
            end
            begin
              @(final_operation[56][6]) ;
            end
            begin
              @(final_operation[56][7]) ;
            end
            begin
              @(final_operation[56][8]) ;
            end
            begin
              @(final_operation[56][9]) ;
            end
            begin
              @(final_operation[56][10]) ;
            end
            begin
              @(final_operation[56][11]) ;
            end
            begin
              @(final_operation[56][12]) ;
            end
            begin
              @(final_operation[56][13]) ;
            end
            begin
              @(final_operation[56][14]) ;
            end
            begin
              @(final_operation[56][15]) ;
            end
            begin
              @(final_operation[56][16]) ;
            end
            begin
              @(final_operation[56][17]) ;
            end
            begin
              @(final_operation[56][18]) ;
            end
            begin
              @(final_operation[56][19]) ;
            end
            begin
              @(final_operation[56][20]) ;
            end
            begin
              @(final_operation[56][21]) ;
            end
            begin
              @(final_operation[56][22]) ;
            end
            begin
              @(final_operation[56][23]) ;
            end
            begin
              @(final_operation[56][24]) ;
            end
            begin
              @(final_operation[56][25]) ;
            end
            begin
              @(final_operation[56][26]) ;
            end
            begin
              @(final_operation[56][27]) ;
            end
            begin
              @(final_operation[56][28]) ;
            end
            begin
              @(final_operation[56][29]) ;
            end
            begin
              @(final_operation[56][30]) ;
            end
            begin
              @(final_operation[56][31]) ;
            end

            begin
              @(final_operation[57][0]) ;
            end
            begin
              @(final_operation[57][1]) ;
            end
            begin
              @(final_operation[57][2]) ;
            end
            begin
              @(final_operation[57][3]) ;
            end
            begin
              @(final_operation[57][4]) ;
            end
            begin
              @(final_operation[57][5]) ;
            end
            begin
              @(final_operation[57][6]) ;
            end
            begin
              @(final_operation[57][7]) ;
            end
            begin
              @(final_operation[57][8]) ;
            end
            begin
              @(final_operation[57][9]) ;
            end
            begin
              @(final_operation[57][10]) ;
            end
            begin
              @(final_operation[57][11]) ;
            end
            begin
              @(final_operation[57][12]) ;
            end
            begin
              @(final_operation[57][13]) ;
            end
            begin
              @(final_operation[57][14]) ;
            end
            begin
              @(final_operation[57][15]) ;
            end
            begin
              @(final_operation[57][16]) ;
            end
            begin
              @(final_operation[57][17]) ;
            end
            begin
              @(final_operation[57][18]) ;
            end
            begin
              @(final_operation[57][19]) ;
            end
            begin
              @(final_operation[57][20]) ;
            end
            begin
              @(final_operation[57][21]) ;
            end
            begin
              @(final_operation[57][22]) ;
            end
            begin
              @(final_operation[57][23]) ;
            end
            begin
              @(final_operation[57][24]) ;
            end
            begin
              @(final_operation[57][25]) ;
            end
            begin
              @(final_operation[57][26]) ;
            end
            begin
              @(final_operation[57][27]) ;
            end
            begin
              @(final_operation[57][28]) ;
            end
            begin
              @(final_operation[57][29]) ;
            end
            begin
              @(final_operation[57][30]) ;
            end
            begin
              @(final_operation[57][31]) ;
            end

            begin
              @(final_operation[58][0]) ;
            end
            begin
              @(final_operation[58][1]) ;
            end
            begin
              @(final_operation[58][2]) ;
            end
            begin
              @(final_operation[58][3]) ;
            end
            begin
              @(final_operation[58][4]) ;
            end
            begin
              @(final_operation[58][5]) ;
            end
            begin
              @(final_operation[58][6]) ;
            end
            begin
              @(final_operation[58][7]) ;
            end
            begin
              @(final_operation[58][8]) ;
            end
            begin
              @(final_operation[58][9]) ;
            end
            begin
              @(final_operation[58][10]) ;
            end
            begin
              @(final_operation[58][11]) ;
            end
            begin
              @(final_operation[58][12]) ;
            end
            begin
              @(final_operation[58][13]) ;
            end
            begin
              @(final_operation[58][14]) ;
            end
            begin
              @(final_operation[58][15]) ;
            end
            begin
              @(final_operation[58][16]) ;
            end
            begin
              @(final_operation[58][17]) ;
            end
            begin
              @(final_operation[58][18]) ;
            end
            begin
              @(final_operation[58][19]) ;
            end
            begin
              @(final_operation[58][20]) ;
            end
            begin
              @(final_operation[58][21]) ;
            end
            begin
              @(final_operation[58][22]) ;
            end
            begin
              @(final_operation[58][23]) ;
            end
            begin
              @(final_operation[58][24]) ;
            end
            begin
              @(final_operation[58][25]) ;
            end
            begin
              @(final_operation[58][26]) ;
            end
            begin
              @(final_operation[58][27]) ;
            end
            begin
              @(final_operation[58][28]) ;
            end
            begin
              @(final_operation[58][29]) ;
            end
            begin
              @(final_operation[58][30]) ;
            end
            begin
              @(final_operation[58][31]) ;
            end

            begin
              @(final_operation[59][0]) ;
            end
            begin
              @(final_operation[59][1]) ;
            end
            begin
              @(final_operation[59][2]) ;
            end
            begin
              @(final_operation[59][3]) ;
            end
            begin
              @(final_operation[59][4]) ;
            end
            begin
              @(final_operation[59][5]) ;
            end
            begin
              @(final_operation[59][6]) ;
            end
            begin
              @(final_operation[59][7]) ;
            end
            begin
              @(final_operation[59][8]) ;
            end
            begin
              @(final_operation[59][9]) ;
            end
            begin
              @(final_operation[59][10]) ;
            end
            begin
              @(final_operation[59][11]) ;
            end
            begin
              @(final_operation[59][12]) ;
            end
            begin
              @(final_operation[59][13]) ;
            end
            begin
              @(final_operation[59][14]) ;
            end
            begin
              @(final_operation[59][15]) ;
            end
            begin
              @(final_operation[59][16]) ;
            end
            begin
              @(final_operation[59][17]) ;
            end
            begin
              @(final_operation[59][18]) ;
            end
            begin
              @(final_operation[59][19]) ;
            end
            begin
              @(final_operation[59][20]) ;
            end
            begin
              @(final_operation[59][21]) ;
            end
            begin
              @(final_operation[59][22]) ;
            end
            begin
              @(final_operation[59][23]) ;
            end
            begin
              @(final_operation[59][24]) ;
            end
            begin
              @(final_operation[59][25]) ;
            end
            begin
              @(final_operation[59][26]) ;
            end
            begin
              @(final_operation[59][27]) ;
            end
            begin
              @(final_operation[59][28]) ;
            end
            begin
              @(final_operation[59][29]) ;
            end
            begin
              @(final_operation[59][30]) ;
            end
            begin
              @(final_operation[59][31]) ;
            end

            begin
              @(final_operation[60][0]) ;
            end
            begin
              @(final_operation[60][1]) ;
            end
            begin
              @(final_operation[60][2]) ;
            end
            begin
              @(final_operation[60][3]) ;
            end
            begin
              @(final_operation[60][4]) ;
            end
            begin
              @(final_operation[60][5]) ;
            end
            begin
              @(final_operation[60][6]) ;
            end
            begin
              @(final_operation[60][7]) ;
            end
            begin
              @(final_operation[60][8]) ;
            end
            begin
              @(final_operation[60][9]) ;
            end
            begin
              @(final_operation[60][10]) ;
            end
            begin
              @(final_operation[60][11]) ;
            end
            begin
              @(final_operation[60][12]) ;
            end
            begin
              @(final_operation[60][13]) ;
            end
            begin
              @(final_operation[60][14]) ;
            end
            begin
              @(final_operation[60][15]) ;
            end
            begin
              @(final_operation[60][16]) ;
            end
            begin
              @(final_operation[60][17]) ;
            end
            begin
              @(final_operation[60][18]) ;
            end
            begin
              @(final_operation[60][19]) ;
            end
            begin
              @(final_operation[60][20]) ;
            end
            begin
              @(final_operation[60][21]) ;
            end
            begin
              @(final_operation[60][22]) ;
            end
            begin
              @(final_operation[60][23]) ;
            end
            begin
              @(final_operation[60][24]) ;
            end
            begin
              @(final_operation[60][25]) ;
            end
            begin
              @(final_operation[60][26]) ;
            end
            begin
              @(final_operation[60][27]) ;
            end
            begin
              @(final_operation[60][28]) ;
            end
            begin
              @(final_operation[60][29]) ;
            end
            begin
              @(final_operation[60][30]) ;
            end
            begin
              @(final_operation[60][31]) ;
            end

            begin
              @(final_operation[61][0]) ;
            end
            begin
              @(final_operation[61][1]) ;
            end
            begin
              @(final_operation[61][2]) ;
            end
            begin
              @(final_operation[61][3]) ;
            end
            begin
              @(final_operation[61][4]) ;
            end
            begin
              @(final_operation[61][5]) ;
            end
            begin
              @(final_operation[61][6]) ;
            end
            begin
              @(final_operation[61][7]) ;
            end
            begin
              @(final_operation[61][8]) ;
            end
            begin
              @(final_operation[61][9]) ;
            end
            begin
              @(final_operation[61][10]) ;
            end
            begin
              @(final_operation[61][11]) ;
            end
            begin
              @(final_operation[61][12]) ;
            end
            begin
              @(final_operation[61][13]) ;
            end
            begin
              @(final_operation[61][14]) ;
            end
            begin
              @(final_operation[61][15]) ;
            end
            begin
              @(final_operation[61][16]) ;
            end
            begin
              @(final_operation[61][17]) ;
            end
            begin
              @(final_operation[61][18]) ;
            end
            begin
              @(final_operation[61][19]) ;
            end
            begin
              @(final_operation[61][20]) ;
            end
            begin
              @(final_operation[61][21]) ;
            end
            begin
              @(final_operation[61][22]) ;
            end
            begin
              @(final_operation[61][23]) ;
            end
            begin
              @(final_operation[61][24]) ;
            end
            begin
              @(final_operation[61][25]) ;
            end
            begin
              @(final_operation[61][26]) ;
            end
            begin
              @(final_operation[61][27]) ;
            end
            begin
              @(final_operation[61][28]) ;
            end
            begin
              @(final_operation[61][29]) ;
            end
            begin
              @(final_operation[61][30]) ;
            end
            begin
              @(final_operation[61][31]) ;
            end

            begin
              @(final_operation[62][0]) ;
            end
            begin
              @(final_operation[62][1]) ;
            end
            begin
              @(final_operation[62][2]) ;
            end
            begin
              @(final_operation[62][3]) ;
            end
            begin
              @(final_operation[62][4]) ;
            end
            begin
              @(final_operation[62][5]) ;
            end
            begin
              @(final_operation[62][6]) ;
            end
            begin
              @(final_operation[62][7]) ;
            end
            begin
              @(final_operation[62][8]) ;
            end
            begin
              @(final_operation[62][9]) ;
            end
            begin
              @(final_operation[62][10]) ;
            end
            begin
              @(final_operation[62][11]) ;
            end
            begin
              @(final_operation[62][12]) ;
            end
            begin
              @(final_operation[62][13]) ;
            end
            begin
              @(final_operation[62][14]) ;
            end
            begin
              @(final_operation[62][15]) ;
            end
            begin
              @(final_operation[62][16]) ;
            end
            begin
              @(final_operation[62][17]) ;
            end
            begin
              @(final_operation[62][18]) ;
            end
            begin
              @(final_operation[62][19]) ;
            end
            begin
              @(final_operation[62][20]) ;
            end
            begin
              @(final_operation[62][21]) ;
            end
            begin
              @(final_operation[62][22]) ;
            end
            begin
              @(final_operation[62][23]) ;
            end
            begin
              @(final_operation[62][24]) ;
            end
            begin
              @(final_operation[62][25]) ;
            end
            begin
              @(final_operation[62][26]) ;
            end
            begin
              @(final_operation[62][27]) ;
            end
            begin
              @(final_operation[62][28]) ;
            end
            begin
              @(final_operation[62][29]) ;
            end
            begin
              @(final_operation[62][30]) ;
            end
            begin
              @(final_operation[62][31]) ;
            end

            begin
              @(final_operation[63][0]) ;
            end
            begin
              @(final_operation[63][1]) ;
            end
            begin
              @(final_operation[63][2]) ;
            end
            begin
              @(final_operation[63][3]) ;
            end
            begin
              @(final_operation[63][4]) ;
            end
            begin
              @(final_operation[63][5]) ;
            end
            begin
              @(final_operation[63][6]) ;
            end
            begin
              @(final_operation[63][7]) ;
            end
            begin
              @(final_operation[63][8]) ;
            end
            begin
              @(final_operation[63][9]) ;
            end
            begin
              @(final_operation[63][10]) ;
            end
            begin
              @(final_operation[63][11]) ;
            end
            begin
              @(final_operation[63][12]) ;
            end
            begin
              @(final_operation[63][13]) ;
            end
            begin
              @(final_operation[63][14]) ;
            end
            begin
              @(final_operation[63][15]) ;
            end
            begin
              @(final_operation[63][16]) ;
            end
            begin
              @(final_operation[63][17]) ;
            end
            begin
              @(final_operation[63][18]) ;
            end
            begin
              @(final_operation[63][19]) ;
            end
            begin
              @(final_operation[63][20]) ;
            end
            begin
              @(final_operation[63][21]) ;
            end
            begin
              @(final_operation[63][22]) ;
            end
            begin
              @(final_operation[63][23]) ;
            end
            begin
              @(final_operation[63][24]) ;
            end
            begin
              @(final_operation[63][25]) ;
            end
            begin
              @(final_operation[63][26]) ;
            end
            begin
              @(final_operation[63][27]) ;
            end
            begin
              @(final_operation[63][28]) ;
            end
            begin
              @(final_operation[63][29]) ;
            end
            begin
              @(final_operation[63][30]) ;
            end
            begin
              @(final_operation[63][31]) ;
            end
