
            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe0__oob_cntl                         ( std__pe0__oob_cntl   ),
            .std__pe0__oob_valid                        ( std__pe0__oob_valid  ),
            .pe0__std__oob_ready                        ( pe0__std__oob_ready  ),
            .std__pe0__oob_type                         ( std__pe0__oob_type   ),
            .std__pe0__oob_data                         ( std__pe0__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe1__oob_cntl                         ( std__pe1__oob_cntl   ),
            .std__pe1__oob_valid                        ( std__pe1__oob_valid  ),
            .pe1__std__oob_ready                        ( pe1__std__oob_ready  ),
            .std__pe1__oob_type                         ( std__pe1__oob_type   ),
            .std__pe1__oob_data                         ( std__pe1__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe2__oob_cntl                         ( std__pe2__oob_cntl   ),
            .std__pe2__oob_valid                        ( std__pe2__oob_valid  ),
            .pe2__std__oob_ready                        ( pe2__std__oob_ready  ),
            .std__pe2__oob_type                         ( std__pe2__oob_type   ),
            .std__pe2__oob_data                         ( std__pe2__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe3__oob_cntl                         ( std__pe3__oob_cntl   ),
            .std__pe3__oob_valid                        ( std__pe3__oob_valid  ),
            .pe3__std__oob_ready                        ( pe3__std__oob_ready  ),
            .std__pe3__oob_type                         ( std__pe3__oob_type   ),
            .std__pe3__oob_data                         ( std__pe3__oob_data   ),

