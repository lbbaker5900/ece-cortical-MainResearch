

            // ##################################################
            // DMA Stream Destination addresses

            // Stream 0 Destination address
            force pe_array_inst.pe_inst[0].pe.lane0_r134 = 32'b000000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane1_r134 = 32'b000000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane2_r134 = 32'b000000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane3_r134 = 32'b000000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane4_r134 = 32'b000000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane5_r134 = 32'b000000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane6_r134 = 32'b000000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane7_r134 = 32'b000000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane8_r134 = 32'b000000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane9_r134 = 32'b000000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane10_r134 = 32'b000000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane11_r134 = 32'b000000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane12_r134 = 32'b000000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane13_r134 = 32'b000000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane14_r134 = 32'b000000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane15_r134 = 32'b000000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane16_r134 = 32'b000000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane17_r134 = 32'b000000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane18_r134 = 32'b000000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane19_r134 = 32'b000000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane20_r134 = 32'b000000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane21_r134 = 32'b000000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane22_r134 = 32'b000000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane23_r134 = 32'b000000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane24_r134 = 32'b000000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane25_r134 = 32'b000000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane26_r134 = 32'b000000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane27_r134 = 32'b000000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane28_r134 = 32'b000000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane29_r134 = 32'b000000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane30_r134 = 32'b000000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.lane31_r134 = 32'b000000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[0].pe.lane0_r135 = 32'b000000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane1_r135 = 32'b000000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane2_r135 = 32'b000000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane3_r135 = 32'b000000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane4_r135 = 32'b000000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane5_r135 = 32'b000000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane6_r135 = 32'b000000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane7_r135 = 32'b000000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane8_r135 = 32'b000000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane9_r135 = 32'b000000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane10_r135 = 32'b000000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane11_r135 = 32'b000000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane12_r135 = 32'b000000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane13_r135 = 32'b000000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane14_r135 = 32'b000000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane15_r135 = 32'b000000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane16_r135 = 32'b000000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane17_r135 = 32'b000000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane18_r135 = 32'b000000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane19_r135 = 32'b000000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane20_r135 = 32'b000000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane21_r135 = 32'b000000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane22_r135 = 32'b000000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane23_r135 = 32'b000000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane24_r135 = 32'b000000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane25_r135 = 32'b000000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane26_r135 = 32'b000000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane27_r135 = 32'b000000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane28_r135 = 32'b000000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane29_r135 = 32'b000000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane30_r135 = 32'b000000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.lane31_r135 = 32'b000000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[1].pe.lane0_r134 = 32'b000001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane1_r134 = 32'b000001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane2_r134 = 32'b000001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane3_r134 = 32'b000001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane4_r134 = 32'b000001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane5_r134 = 32'b000001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane6_r134 = 32'b000001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane7_r134 = 32'b000001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane8_r134 = 32'b000001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane9_r134 = 32'b000001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane10_r134 = 32'b000001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane11_r134 = 32'b000001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane12_r134 = 32'b000001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane13_r134 = 32'b000001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane14_r134 = 32'b000001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane15_r134 = 32'b000001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane16_r134 = 32'b000001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane17_r134 = 32'b000001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane18_r134 = 32'b000001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane19_r134 = 32'b000001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane20_r134 = 32'b000001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane21_r134 = 32'b000001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane22_r134 = 32'b000001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane23_r134 = 32'b000001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane24_r134 = 32'b000001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane25_r134 = 32'b000001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane26_r134 = 32'b000001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane27_r134 = 32'b000001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane28_r134 = 32'b000001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane29_r134 = 32'b000001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane30_r134 = 32'b000001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.lane31_r134 = 32'b000001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[1].pe.lane0_r135 = 32'b000001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane1_r135 = 32'b000001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane2_r135 = 32'b000001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane3_r135 = 32'b000001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane4_r135 = 32'b000001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane5_r135 = 32'b000001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane6_r135 = 32'b000001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane7_r135 = 32'b000001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane8_r135 = 32'b000001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane9_r135 = 32'b000001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane10_r135 = 32'b000001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane11_r135 = 32'b000001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane12_r135 = 32'b000001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane13_r135 = 32'b000001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane14_r135 = 32'b000001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane15_r135 = 32'b000001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane16_r135 = 32'b000001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane17_r135 = 32'b000001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane18_r135 = 32'b000001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane19_r135 = 32'b000001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane20_r135 = 32'b000001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane21_r135 = 32'b000001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane22_r135 = 32'b000001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane23_r135 = 32'b000001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane24_r135 = 32'b000001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane25_r135 = 32'b000001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane26_r135 = 32'b000001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane27_r135 = 32'b000001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane28_r135 = 32'b000001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane29_r135 = 32'b000001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane30_r135 = 32'b000001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.lane31_r135 = 32'b000001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[2].pe.lane0_r134 = 32'b000010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane1_r134 = 32'b000010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane2_r134 = 32'b000010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane3_r134 = 32'b000010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane4_r134 = 32'b000010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane5_r134 = 32'b000010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane6_r134 = 32'b000010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane7_r134 = 32'b000010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane8_r134 = 32'b000010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane9_r134 = 32'b000010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane10_r134 = 32'b000010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane11_r134 = 32'b000010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane12_r134 = 32'b000010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane13_r134 = 32'b000010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane14_r134 = 32'b000010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane15_r134 = 32'b000010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane16_r134 = 32'b000010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane17_r134 = 32'b000010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane18_r134 = 32'b000010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane19_r134 = 32'b000010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane20_r134 = 32'b000010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane21_r134 = 32'b000010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane22_r134 = 32'b000010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane23_r134 = 32'b000010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane24_r134 = 32'b000010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane25_r134 = 32'b000010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane26_r134 = 32'b000010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane27_r134 = 32'b000010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane28_r134 = 32'b000010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane29_r134 = 32'b000010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane30_r134 = 32'b000010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.lane31_r134 = 32'b000010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[2].pe.lane0_r135 = 32'b000010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane1_r135 = 32'b000010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane2_r135 = 32'b000010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane3_r135 = 32'b000010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane4_r135 = 32'b000010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane5_r135 = 32'b000010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane6_r135 = 32'b000010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane7_r135 = 32'b000010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane8_r135 = 32'b000010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane9_r135 = 32'b000010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane10_r135 = 32'b000010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane11_r135 = 32'b000010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane12_r135 = 32'b000010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane13_r135 = 32'b000010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane14_r135 = 32'b000010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane15_r135 = 32'b000010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane16_r135 = 32'b000010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane17_r135 = 32'b000010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane18_r135 = 32'b000010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane19_r135 = 32'b000010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane20_r135 = 32'b000010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane21_r135 = 32'b000010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane22_r135 = 32'b000010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane23_r135 = 32'b000010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane24_r135 = 32'b000010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane25_r135 = 32'b000010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane26_r135 = 32'b000010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane27_r135 = 32'b000010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane28_r135 = 32'b000010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane29_r135 = 32'b000010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane30_r135 = 32'b000010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.lane31_r135 = 32'b000010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[3].pe.lane0_r134 = 32'b000011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane1_r134 = 32'b000011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane2_r134 = 32'b000011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane3_r134 = 32'b000011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane4_r134 = 32'b000011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane5_r134 = 32'b000011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane6_r134 = 32'b000011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane7_r134 = 32'b000011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane8_r134 = 32'b000011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane9_r134 = 32'b000011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane10_r134 = 32'b000011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane11_r134 = 32'b000011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane12_r134 = 32'b000011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane13_r134 = 32'b000011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane14_r134 = 32'b000011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane15_r134 = 32'b000011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane16_r134 = 32'b000011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane17_r134 = 32'b000011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane18_r134 = 32'b000011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane19_r134 = 32'b000011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane20_r134 = 32'b000011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane21_r134 = 32'b000011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane22_r134 = 32'b000011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane23_r134 = 32'b000011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane24_r134 = 32'b000011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane25_r134 = 32'b000011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane26_r134 = 32'b000011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane27_r134 = 32'b000011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane28_r134 = 32'b000011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane29_r134 = 32'b000011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane30_r134 = 32'b000011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.lane31_r134 = 32'b000011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[3].pe.lane0_r135 = 32'b000011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane1_r135 = 32'b000011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane2_r135 = 32'b000011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane3_r135 = 32'b000011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane4_r135 = 32'b000011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane5_r135 = 32'b000011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane6_r135 = 32'b000011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane7_r135 = 32'b000011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane8_r135 = 32'b000011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane9_r135 = 32'b000011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane10_r135 = 32'b000011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane11_r135 = 32'b000011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane12_r135 = 32'b000011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane13_r135 = 32'b000011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane14_r135 = 32'b000011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane15_r135 = 32'b000011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane16_r135 = 32'b000011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane17_r135 = 32'b000011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane18_r135 = 32'b000011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane19_r135 = 32'b000011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane20_r135 = 32'b000011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane21_r135 = 32'b000011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane22_r135 = 32'b000011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane23_r135 = 32'b000011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane24_r135 = 32'b000011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane25_r135 = 32'b000011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane26_r135 = 32'b000011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane27_r135 = 32'b000011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane28_r135 = 32'b000011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane29_r135 = 32'b000011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane30_r135 = 32'b000011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.lane31_r135 = 32'b000011_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[4].pe.lane0_r134 = 32'b000100_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane1_r134 = 32'b000100_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane2_r134 = 32'b000100_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane3_r134 = 32'b000100_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane4_r134 = 32'b000100_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane5_r134 = 32'b000100_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane6_r134 = 32'b000100_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane7_r134 = 32'b000100_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane8_r134 = 32'b000100_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane9_r134 = 32'b000100_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane10_r134 = 32'b000100_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane11_r134 = 32'b000100_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane12_r134 = 32'b000100_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane13_r134 = 32'b000100_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane14_r134 = 32'b000100_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane15_r134 = 32'b000100_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane16_r134 = 32'b000100_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane17_r134 = 32'b000100_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane18_r134 = 32'b000100_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane19_r134 = 32'b000100_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane20_r134 = 32'b000100_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane21_r134 = 32'b000100_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane22_r134 = 32'b000100_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane23_r134 = 32'b000100_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane24_r134 = 32'b000100_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane25_r134 = 32'b000100_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane26_r134 = 32'b000100_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane27_r134 = 32'b000100_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane28_r134 = 32'b000100_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane29_r134 = 32'b000100_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane30_r134 = 32'b000100_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.lane31_r134 = 32'b000100_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[4].pe.lane0_r135 = 32'b000100_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane1_r135 = 32'b000100_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane2_r135 = 32'b000100_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane3_r135 = 32'b000100_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane4_r135 = 32'b000100_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane5_r135 = 32'b000100_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane6_r135 = 32'b000100_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane7_r135 = 32'b000100_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane8_r135 = 32'b000100_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane9_r135 = 32'b000100_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane10_r135 = 32'b000100_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane11_r135 = 32'b000100_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane12_r135 = 32'b000100_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane13_r135 = 32'b000100_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane14_r135 = 32'b000100_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane15_r135 = 32'b000100_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane16_r135 = 32'b000100_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane17_r135 = 32'b000100_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane18_r135 = 32'b000100_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane19_r135 = 32'b000100_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane20_r135 = 32'b000100_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane21_r135 = 32'b000100_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane22_r135 = 32'b000100_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane23_r135 = 32'b000100_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane24_r135 = 32'b000100_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane25_r135 = 32'b000100_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane26_r135 = 32'b000100_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane27_r135 = 32'b000100_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane28_r135 = 32'b000100_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane29_r135 = 32'b000100_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane30_r135 = 32'b000100_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.lane31_r135 = 32'b000100_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[5].pe.lane0_r134 = 32'b000101_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane1_r134 = 32'b000101_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane2_r134 = 32'b000101_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane3_r134 = 32'b000101_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane4_r134 = 32'b000101_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane5_r134 = 32'b000101_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane6_r134 = 32'b000101_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane7_r134 = 32'b000101_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane8_r134 = 32'b000101_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane9_r134 = 32'b000101_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane10_r134 = 32'b000101_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane11_r134 = 32'b000101_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane12_r134 = 32'b000101_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane13_r134 = 32'b000101_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane14_r134 = 32'b000101_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane15_r134 = 32'b000101_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane16_r134 = 32'b000101_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane17_r134 = 32'b000101_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane18_r134 = 32'b000101_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane19_r134 = 32'b000101_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane20_r134 = 32'b000101_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane21_r134 = 32'b000101_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane22_r134 = 32'b000101_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane23_r134 = 32'b000101_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane24_r134 = 32'b000101_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane25_r134 = 32'b000101_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane26_r134 = 32'b000101_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane27_r134 = 32'b000101_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane28_r134 = 32'b000101_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane29_r134 = 32'b000101_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane30_r134 = 32'b000101_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.lane31_r134 = 32'b000101_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[5].pe.lane0_r135 = 32'b000101_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane1_r135 = 32'b000101_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane2_r135 = 32'b000101_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane3_r135 = 32'b000101_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane4_r135 = 32'b000101_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane5_r135 = 32'b000101_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane6_r135 = 32'b000101_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane7_r135 = 32'b000101_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane8_r135 = 32'b000101_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane9_r135 = 32'b000101_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane10_r135 = 32'b000101_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane11_r135 = 32'b000101_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane12_r135 = 32'b000101_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane13_r135 = 32'b000101_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane14_r135 = 32'b000101_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane15_r135 = 32'b000101_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane16_r135 = 32'b000101_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane17_r135 = 32'b000101_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane18_r135 = 32'b000101_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane19_r135 = 32'b000101_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane20_r135 = 32'b000101_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane21_r135 = 32'b000101_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane22_r135 = 32'b000101_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane23_r135 = 32'b000101_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane24_r135 = 32'b000101_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane25_r135 = 32'b000101_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane26_r135 = 32'b000101_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane27_r135 = 32'b000101_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane28_r135 = 32'b000101_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane29_r135 = 32'b000101_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane30_r135 = 32'b000101_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.lane31_r135 = 32'b000101_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[6].pe.lane0_r134 = 32'b000110_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane1_r134 = 32'b000110_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane2_r134 = 32'b000110_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane3_r134 = 32'b000110_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane4_r134 = 32'b000110_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane5_r134 = 32'b000110_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane6_r134 = 32'b000110_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane7_r134 = 32'b000110_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane8_r134 = 32'b000110_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane9_r134 = 32'b000110_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane10_r134 = 32'b000110_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane11_r134 = 32'b000110_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane12_r134 = 32'b000110_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane13_r134 = 32'b000110_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane14_r134 = 32'b000110_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane15_r134 = 32'b000110_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane16_r134 = 32'b000110_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane17_r134 = 32'b000110_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane18_r134 = 32'b000110_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane19_r134 = 32'b000110_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane20_r134 = 32'b000110_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane21_r134 = 32'b000110_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane22_r134 = 32'b000110_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane23_r134 = 32'b000110_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane24_r134 = 32'b000110_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane25_r134 = 32'b000110_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane26_r134 = 32'b000110_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane27_r134 = 32'b000110_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane28_r134 = 32'b000110_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane29_r134 = 32'b000110_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane30_r134 = 32'b000110_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.lane31_r134 = 32'b000110_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[6].pe.lane0_r135 = 32'b000110_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane1_r135 = 32'b000110_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane2_r135 = 32'b000110_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane3_r135 = 32'b000110_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane4_r135 = 32'b000110_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane5_r135 = 32'b000110_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane6_r135 = 32'b000110_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane7_r135 = 32'b000110_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane8_r135 = 32'b000110_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane9_r135 = 32'b000110_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane10_r135 = 32'b000110_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane11_r135 = 32'b000110_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane12_r135 = 32'b000110_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane13_r135 = 32'b000110_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane14_r135 = 32'b000110_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane15_r135 = 32'b000110_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane16_r135 = 32'b000110_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane17_r135 = 32'b000110_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane18_r135 = 32'b000110_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane19_r135 = 32'b000110_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane20_r135 = 32'b000110_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane21_r135 = 32'b000110_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane22_r135 = 32'b000110_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane23_r135 = 32'b000110_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane24_r135 = 32'b000110_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane25_r135 = 32'b000110_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane26_r135 = 32'b000110_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane27_r135 = 32'b000110_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane28_r135 = 32'b000110_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane29_r135 = 32'b000110_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane30_r135 = 32'b000110_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.lane31_r135 = 32'b000110_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[7].pe.lane0_r134 = 32'b000111_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane1_r134 = 32'b000111_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane2_r134 = 32'b000111_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane3_r134 = 32'b000111_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane4_r134 = 32'b000111_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane5_r134 = 32'b000111_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane6_r134 = 32'b000111_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane7_r134 = 32'b000111_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane8_r134 = 32'b000111_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane9_r134 = 32'b000111_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane10_r134 = 32'b000111_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane11_r134 = 32'b000111_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane12_r134 = 32'b000111_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane13_r134 = 32'b000111_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane14_r134 = 32'b000111_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane15_r134 = 32'b000111_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane16_r134 = 32'b000111_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane17_r134 = 32'b000111_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane18_r134 = 32'b000111_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane19_r134 = 32'b000111_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane20_r134 = 32'b000111_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane21_r134 = 32'b000111_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane22_r134 = 32'b000111_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane23_r134 = 32'b000111_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane24_r134 = 32'b000111_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane25_r134 = 32'b000111_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane26_r134 = 32'b000111_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane27_r134 = 32'b000111_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane28_r134 = 32'b000111_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane29_r134 = 32'b000111_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane30_r134 = 32'b000111_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.lane31_r134 = 32'b000111_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[7].pe.lane0_r135 = 32'b000111_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane1_r135 = 32'b000111_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane2_r135 = 32'b000111_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane3_r135 = 32'b000111_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane4_r135 = 32'b000111_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane5_r135 = 32'b000111_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane6_r135 = 32'b000111_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane7_r135 = 32'b000111_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane8_r135 = 32'b000111_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane9_r135 = 32'b000111_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane10_r135 = 32'b000111_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane11_r135 = 32'b000111_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane12_r135 = 32'b000111_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane13_r135 = 32'b000111_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane14_r135 = 32'b000111_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane15_r135 = 32'b000111_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane16_r135 = 32'b000111_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane17_r135 = 32'b000111_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane18_r135 = 32'b000111_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane19_r135 = 32'b000111_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane20_r135 = 32'b000111_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane21_r135 = 32'b000111_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane22_r135 = 32'b000111_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane23_r135 = 32'b000111_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane24_r135 = 32'b000111_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane25_r135 = 32'b000111_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane26_r135 = 32'b000111_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane27_r135 = 32'b000111_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane28_r135 = 32'b000111_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane29_r135 = 32'b000111_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane30_r135 = 32'b000111_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.lane31_r135 = 32'b000111_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[8].pe.lane0_r134 = 32'b001000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane1_r134 = 32'b001000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane2_r134 = 32'b001000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane3_r134 = 32'b001000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane4_r134 = 32'b001000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane5_r134 = 32'b001000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane6_r134 = 32'b001000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane7_r134 = 32'b001000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane8_r134 = 32'b001000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane9_r134 = 32'b001000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane10_r134 = 32'b001000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane11_r134 = 32'b001000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane12_r134 = 32'b001000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane13_r134 = 32'b001000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane14_r134 = 32'b001000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane15_r134 = 32'b001000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane16_r134 = 32'b001000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane17_r134 = 32'b001000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane18_r134 = 32'b001000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane19_r134 = 32'b001000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane20_r134 = 32'b001000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane21_r134 = 32'b001000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane22_r134 = 32'b001000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane23_r134 = 32'b001000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane24_r134 = 32'b001000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane25_r134 = 32'b001000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane26_r134 = 32'b001000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane27_r134 = 32'b001000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane28_r134 = 32'b001000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane29_r134 = 32'b001000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane30_r134 = 32'b001000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.lane31_r134 = 32'b001000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[8].pe.lane0_r135 = 32'b001000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane1_r135 = 32'b001000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane2_r135 = 32'b001000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane3_r135 = 32'b001000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane4_r135 = 32'b001000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane5_r135 = 32'b001000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane6_r135 = 32'b001000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane7_r135 = 32'b001000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane8_r135 = 32'b001000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane9_r135 = 32'b001000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane10_r135 = 32'b001000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane11_r135 = 32'b001000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane12_r135 = 32'b001000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane13_r135 = 32'b001000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane14_r135 = 32'b001000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane15_r135 = 32'b001000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane16_r135 = 32'b001000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane17_r135 = 32'b001000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane18_r135 = 32'b001000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane19_r135 = 32'b001000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane20_r135 = 32'b001000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane21_r135 = 32'b001000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane22_r135 = 32'b001000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane23_r135 = 32'b001000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane24_r135 = 32'b001000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane25_r135 = 32'b001000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane26_r135 = 32'b001000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane27_r135 = 32'b001000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane28_r135 = 32'b001000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane29_r135 = 32'b001000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane30_r135 = 32'b001000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.lane31_r135 = 32'b001000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[9].pe.lane0_r134 = 32'b001001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane1_r134 = 32'b001001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane2_r134 = 32'b001001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane3_r134 = 32'b001001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane4_r134 = 32'b001001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane5_r134 = 32'b001001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane6_r134 = 32'b001001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane7_r134 = 32'b001001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane8_r134 = 32'b001001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane9_r134 = 32'b001001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane10_r134 = 32'b001001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane11_r134 = 32'b001001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane12_r134 = 32'b001001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane13_r134 = 32'b001001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane14_r134 = 32'b001001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane15_r134 = 32'b001001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane16_r134 = 32'b001001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane17_r134 = 32'b001001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane18_r134 = 32'b001001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane19_r134 = 32'b001001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane20_r134 = 32'b001001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane21_r134 = 32'b001001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane22_r134 = 32'b001001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane23_r134 = 32'b001001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane24_r134 = 32'b001001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane25_r134 = 32'b001001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane26_r134 = 32'b001001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane27_r134 = 32'b001001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane28_r134 = 32'b001001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane29_r134 = 32'b001001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane30_r134 = 32'b001001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.lane31_r134 = 32'b001001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[9].pe.lane0_r135 = 32'b001001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane1_r135 = 32'b001001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane2_r135 = 32'b001001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane3_r135 = 32'b001001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane4_r135 = 32'b001001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane5_r135 = 32'b001001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane6_r135 = 32'b001001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane7_r135 = 32'b001001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane8_r135 = 32'b001001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane9_r135 = 32'b001001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane10_r135 = 32'b001001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane11_r135 = 32'b001001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane12_r135 = 32'b001001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane13_r135 = 32'b001001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane14_r135 = 32'b001001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane15_r135 = 32'b001001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane16_r135 = 32'b001001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane17_r135 = 32'b001001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane18_r135 = 32'b001001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane19_r135 = 32'b001001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane20_r135 = 32'b001001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane21_r135 = 32'b001001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane22_r135 = 32'b001001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane23_r135 = 32'b001001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane24_r135 = 32'b001001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane25_r135 = 32'b001001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane26_r135 = 32'b001001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane27_r135 = 32'b001001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane28_r135 = 32'b001001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane29_r135 = 32'b001001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane30_r135 = 32'b001001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.lane31_r135 = 32'b001001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[10].pe.lane0_r134 = 32'b001010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane1_r134 = 32'b001010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane2_r134 = 32'b001010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane3_r134 = 32'b001010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane4_r134 = 32'b001010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane5_r134 = 32'b001010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane6_r134 = 32'b001010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane7_r134 = 32'b001010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane8_r134 = 32'b001010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane9_r134 = 32'b001010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane10_r134 = 32'b001010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane11_r134 = 32'b001010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane12_r134 = 32'b001010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane13_r134 = 32'b001010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane14_r134 = 32'b001010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane15_r134 = 32'b001010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane16_r134 = 32'b001010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane17_r134 = 32'b001010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane18_r134 = 32'b001010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane19_r134 = 32'b001010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane20_r134 = 32'b001010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane21_r134 = 32'b001010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane22_r134 = 32'b001010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane23_r134 = 32'b001010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane24_r134 = 32'b001010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane25_r134 = 32'b001010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane26_r134 = 32'b001010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane27_r134 = 32'b001010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane28_r134 = 32'b001010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane29_r134 = 32'b001010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane30_r134 = 32'b001010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.lane31_r134 = 32'b001010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[10].pe.lane0_r135 = 32'b001010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane1_r135 = 32'b001010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane2_r135 = 32'b001010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane3_r135 = 32'b001010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane4_r135 = 32'b001010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane5_r135 = 32'b001010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane6_r135 = 32'b001010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane7_r135 = 32'b001010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane8_r135 = 32'b001010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane9_r135 = 32'b001010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane10_r135 = 32'b001010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane11_r135 = 32'b001010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane12_r135 = 32'b001010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane13_r135 = 32'b001010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane14_r135 = 32'b001010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane15_r135 = 32'b001010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane16_r135 = 32'b001010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane17_r135 = 32'b001010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane18_r135 = 32'b001010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane19_r135 = 32'b001010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane20_r135 = 32'b001010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane21_r135 = 32'b001010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane22_r135 = 32'b001010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane23_r135 = 32'b001010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane24_r135 = 32'b001010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane25_r135 = 32'b001010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane26_r135 = 32'b001010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane27_r135 = 32'b001010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane28_r135 = 32'b001010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane29_r135 = 32'b001010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane30_r135 = 32'b001010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.lane31_r135 = 32'b001010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[11].pe.lane0_r134 = 32'b001011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane1_r134 = 32'b001011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane2_r134 = 32'b001011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane3_r134 = 32'b001011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane4_r134 = 32'b001011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane5_r134 = 32'b001011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane6_r134 = 32'b001011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane7_r134 = 32'b001011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane8_r134 = 32'b001011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane9_r134 = 32'b001011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane10_r134 = 32'b001011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane11_r134 = 32'b001011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane12_r134 = 32'b001011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane13_r134 = 32'b001011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane14_r134 = 32'b001011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane15_r134 = 32'b001011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane16_r134 = 32'b001011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane17_r134 = 32'b001011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane18_r134 = 32'b001011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane19_r134 = 32'b001011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane20_r134 = 32'b001011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane21_r134 = 32'b001011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane22_r134 = 32'b001011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane23_r134 = 32'b001011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane24_r134 = 32'b001011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane25_r134 = 32'b001011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane26_r134 = 32'b001011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane27_r134 = 32'b001011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane28_r134 = 32'b001011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane29_r134 = 32'b001011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane30_r134 = 32'b001011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.lane31_r134 = 32'b001011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[11].pe.lane0_r135 = 32'b001011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane1_r135 = 32'b001011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane2_r135 = 32'b001011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane3_r135 = 32'b001011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane4_r135 = 32'b001011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane5_r135 = 32'b001011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane6_r135 = 32'b001011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane7_r135 = 32'b001011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane8_r135 = 32'b001011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane9_r135 = 32'b001011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane10_r135 = 32'b001011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane11_r135 = 32'b001011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane12_r135 = 32'b001011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane13_r135 = 32'b001011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane14_r135 = 32'b001011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane15_r135 = 32'b001011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane16_r135 = 32'b001011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane17_r135 = 32'b001011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane18_r135 = 32'b001011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane19_r135 = 32'b001011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane20_r135 = 32'b001011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane21_r135 = 32'b001011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane22_r135 = 32'b001011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane23_r135 = 32'b001011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane24_r135 = 32'b001011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane25_r135 = 32'b001011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane26_r135 = 32'b001011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane27_r135 = 32'b001011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane28_r135 = 32'b001011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane29_r135 = 32'b001011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane30_r135 = 32'b001011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.lane31_r135 = 32'b001011_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[12].pe.lane0_r134 = 32'b001100_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane1_r134 = 32'b001100_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane2_r134 = 32'b001100_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane3_r134 = 32'b001100_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane4_r134 = 32'b001100_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane5_r134 = 32'b001100_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane6_r134 = 32'b001100_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane7_r134 = 32'b001100_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane8_r134 = 32'b001100_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane9_r134 = 32'b001100_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane10_r134 = 32'b001100_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane11_r134 = 32'b001100_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane12_r134 = 32'b001100_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane13_r134 = 32'b001100_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane14_r134 = 32'b001100_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane15_r134 = 32'b001100_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane16_r134 = 32'b001100_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane17_r134 = 32'b001100_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane18_r134 = 32'b001100_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane19_r134 = 32'b001100_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane20_r134 = 32'b001100_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane21_r134 = 32'b001100_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane22_r134 = 32'b001100_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane23_r134 = 32'b001100_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane24_r134 = 32'b001100_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane25_r134 = 32'b001100_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane26_r134 = 32'b001100_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane27_r134 = 32'b001100_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane28_r134 = 32'b001100_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane29_r134 = 32'b001100_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane30_r134 = 32'b001100_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.lane31_r134 = 32'b001100_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[12].pe.lane0_r135 = 32'b001100_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane1_r135 = 32'b001100_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane2_r135 = 32'b001100_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane3_r135 = 32'b001100_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane4_r135 = 32'b001100_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane5_r135 = 32'b001100_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane6_r135 = 32'b001100_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane7_r135 = 32'b001100_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane8_r135 = 32'b001100_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane9_r135 = 32'b001100_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane10_r135 = 32'b001100_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane11_r135 = 32'b001100_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane12_r135 = 32'b001100_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane13_r135 = 32'b001100_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane14_r135 = 32'b001100_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane15_r135 = 32'b001100_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane16_r135 = 32'b001100_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane17_r135 = 32'b001100_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane18_r135 = 32'b001100_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane19_r135 = 32'b001100_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane20_r135 = 32'b001100_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane21_r135 = 32'b001100_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane22_r135 = 32'b001100_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane23_r135 = 32'b001100_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane24_r135 = 32'b001100_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane25_r135 = 32'b001100_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane26_r135 = 32'b001100_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane27_r135 = 32'b001100_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane28_r135 = 32'b001100_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane29_r135 = 32'b001100_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane30_r135 = 32'b001100_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.lane31_r135 = 32'b001100_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[13].pe.lane0_r134 = 32'b001101_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane1_r134 = 32'b001101_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane2_r134 = 32'b001101_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane3_r134 = 32'b001101_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane4_r134 = 32'b001101_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane5_r134 = 32'b001101_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane6_r134 = 32'b001101_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane7_r134 = 32'b001101_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane8_r134 = 32'b001101_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane9_r134 = 32'b001101_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane10_r134 = 32'b001101_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane11_r134 = 32'b001101_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane12_r134 = 32'b001101_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane13_r134 = 32'b001101_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane14_r134 = 32'b001101_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane15_r134 = 32'b001101_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane16_r134 = 32'b001101_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane17_r134 = 32'b001101_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane18_r134 = 32'b001101_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane19_r134 = 32'b001101_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane20_r134 = 32'b001101_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane21_r134 = 32'b001101_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane22_r134 = 32'b001101_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane23_r134 = 32'b001101_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane24_r134 = 32'b001101_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane25_r134 = 32'b001101_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane26_r134 = 32'b001101_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane27_r134 = 32'b001101_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane28_r134 = 32'b001101_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane29_r134 = 32'b001101_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane30_r134 = 32'b001101_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.lane31_r134 = 32'b001101_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[13].pe.lane0_r135 = 32'b001101_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane1_r135 = 32'b001101_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane2_r135 = 32'b001101_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane3_r135 = 32'b001101_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane4_r135 = 32'b001101_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane5_r135 = 32'b001101_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane6_r135 = 32'b001101_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane7_r135 = 32'b001101_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane8_r135 = 32'b001101_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane9_r135 = 32'b001101_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane10_r135 = 32'b001101_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane11_r135 = 32'b001101_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane12_r135 = 32'b001101_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane13_r135 = 32'b001101_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane14_r135 = 32'b001101_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane15_r135 = 32'b001101_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane16_r135 = 32'b001101_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane17_r135 = 32'b001101_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane18_r135 = 32'b001101_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane19_r135 = 32'b001101_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane20_r135 = 32'b001101_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane21_r135 = 32'b001101_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane22_r135 = 32'b001101_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane23_r135 = 32'b001101_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane24_r135 = 32'b001101_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane25_r135 = 32'b001101_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane26_r135 = 32'b001101_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane27_r135 = 32'b001101_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane28_r135 = 32'b001101_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane29_r135 = 32'b001101_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane30_r135 = 32'b001101_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.lane31_r135 = 32'b001101_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[14].pe.lane0_r134 = 32'b001110_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane1_r134 = 32'b001110_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane2_r134 = 32'b001110_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane3_r134 = 32'b001110_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane4_r134 = 32'b001110_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane5_r134 = 32'b001110_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane6_r134 = 32'b001110_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane7_r134 = 32'b001110_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane8_r134 = 32'b001110_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane9_r134 = 32'b001110_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane10_r134 = 32'b001110_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane11_r134 = 32'b001110_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane12_r134 = 32'b001110_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane13_r134 = 32'b001110_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane14_r134 = 32'b001110_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane15_r134 = 32'b001110_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane16_r134 = 32'b001110_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane17_r134 = 32'b001110_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane18_r134 = 32'b001110_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane19_r134 = 32'b001110_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane20_r134 = 32'b001110_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane21_r134 = 32'b001110_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane22_r134 = 32'b001110_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane23_r134 = 32'b001110_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane24_r134 = 32'b001110_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane25_r134 = 32'b001110_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane26_r134 = 32'b001110_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane27_r134 = 32'b001110_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane28_r134 = 32'b001110_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane29_r134 = 32'b001110_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane30_r134 = 32'b001110_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.lane31_r134 = 32'b001110_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[14].pe.lane0_r135 = 32'b001110_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane1_r135 = 32'b001110_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane2_r135 = 32'b001110_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane3_r135 = 32'b001110_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane4_r135 = 32'b001110_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane5_r135 = 32'b001110_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane6_r135 = 32'b001110_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane7_r135 = 32'b001110_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane8_r135 = 32'b001110_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane9_r135 = 32'b001110_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane10_r135 = 32'b001110_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane11_r135 = 32'b001110_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane12_r135 = 32'b001110_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane13_r135 = 32'b001110_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane14_r135 = 32'b001110_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane15_r135 = 32'b001110_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane16_r135 = 32'b001110_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane17_r135 = 32'b001110_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane18_r135 = 32'b001110_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane19_r135 = 32'b001110_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane20_r135 = 32'b001110_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane21_r135 = 32'b001110_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane22_r135 = 32'b001110_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane23_r135 = 32'b001110_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane24_r135 = 32'b001110_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane25_r135 = 32'b001110_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane26_r135 = 32'b001110_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane27_r135 = 32'b001110_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane28_r135 = 32'b001110_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane29_r135 = 32'b001110_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane30_r135 = 32'b001110_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.lane31_r135 = 32'b001110_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[15].pe.lane0_r134 = 32'b001111_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane1_r134 = 32'b001111_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane2_r134 = 32'b001111_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane3_r134 = 32'b001111_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane4_r134 = 32'b001111_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane5_r134 = 32'b001111_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane6_r134 = 32'b001111_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane7_r134 = 32'b001111_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane8_r134 = 32'b001111_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane9_r134 = 32'b001111_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane10_r134 = 32'b001111_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane11_r134 = 32'b001111_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane12_r134 = 32'b001111_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane13_r134 = 32'b001111_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane14_r134 = 32'b001111_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane15_r134 = 32'b001111_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane16_r134 = 32'b001111_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane17_r134 = 32'b001111_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane18_r134 = 32'b001111_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane19_r134 = 32'b001111_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane20_r134 = 32'b001111_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane21_r134 = 32'b001111_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane22_r134 = 32'b001111_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane23_r134 = 32'b001111_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane24_r134 = 32'b001111_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane25_r134 = 32'b001111_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane26_r134 = 32'b001111_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane27_r134 = 32'b001111_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane28_r134 = 32'b001111_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane29_r134 = 32'b001111_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane30_r134 = 32'b001111_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.lane31_r134 = 32'b001111_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[15].pe.lane0_r135 = 32'b001111_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane1_r135 = 32'b001111_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane2_r135 = 32'b001111_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane3_r135 = 32'b001111_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane4_r135 = 32'b001111_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane5_r135 = 32'b001111_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane6_r135 = 32'b001111_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane7_r135 = 32'b001111_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane8_r135 = 32'b001111_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane9_r135 = 32'b001111_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane10_r135 = 32'b001111_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane11_r135 = 32'b001111_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane12_r135 = 32'b001111_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane13_r135 = 32'b001111_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane14_r135 = 32'b001111_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane15_r135 = 32'b001111_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane16_r135 = 32'b001111_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane17_r135 = 32'b001111_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane18_r135 = 32'b001111_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane19_r135 = 32'b001111_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane20_r135 = 32'b001111_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane21_r135 = 32'b001111_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane22_r135 = 32'b001111_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane23_r135 = 32'b001111_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane24_r135 = 32'b001111_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane25_r135 = 32'b001111_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane26_r135 = 32'b001111_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane27_r135 = 32'b001111_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane28_r135 = 32'b001111_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane29_r135 = 32'b001111_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane30_r135 = 32'b001111_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.lane31_r135 = 32'b001111_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[16].pe.lane0_r134 = 32'b010000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane1_r134 = 32'b010000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane2_r134 = 32'b010000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane3_r134 = 32'b010000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane4_r134 = 32'b010000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane5_r134 = 32'b010000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane6_r134 = 32'b010000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane7_r134 = 32'b010000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane8_r134 = 32'b010000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane9_r134 = 32'b010000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane10_r134 = 32'b010000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane11_r134 = 32'b010000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane12_r134 = 32'b010000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane13_r134 = 32'b010000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane14_r134 = 32'b010000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane15_r134 = 32'b010000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane16_r134 = 32'b010000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane17_r134 = 32'b010000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane18_r134 = 32'b010000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane19_r134 = 32'b010000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane20_r134 = 32'b010000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane21_r134 = 32'b010000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane22_r134 = 32'b010000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane23_r134 = 32'b010000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane24_r134 = 32'b010000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane25_r134 = 32'b010000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane26_r134 = 32'b010000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane27_r134 = 32'b010000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane28_r134 = 32'b010000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane29_r134 = 32'b010000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane30_r134 = 32'b010000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.lane31_r134 = 32'b010000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[16].pe.lane0_r135 = 32'b010000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane1_r135 = 32'b010000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane2_r135 = 32'b010000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane3_r135 = 32'b010000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane4_r135 = 32'b010000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane5_r135 = 32'b010000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane6_r135 = 32'b010000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane7_r135 = 32'b010000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane8_r135 = 32'b010000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane9_r135 = 32'b010000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane10_r135 = 32'b010000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane11_r135 = 32'b010000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane12_r135 = 32'b010000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane13_r135 = 32'b010000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane14_r135 = 32'b010000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane15_r135 = 32'b010000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane16_r135 = 32'b010000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane17_r135 = 32'b010000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane18_r135 = 32'b010000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane19_r135 = 32'b010000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane20_r135 = 32'b010000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane21_r135 = 32'b010000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane22_r135 = 32'b010000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane23_r135 = 32'b010000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane24_r135 = 32'b010000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane25_r135 = 32'b010000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane26_r135 = 32'b010000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane27_r135 = 32'b010000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane28_r135 = 32'b010000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane29_r135 = 32'b010000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane30_r135 = 32'b010000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.lane31_r135 = 32'b010000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[17].pe.lane0_r134 = 32'b010001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane1_r134 = 32'b010001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane2_r134 = 32'b010001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane3_r134 = 32'b010001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane4_r134 = 32'b010001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane5_r134 = 32'b010001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane6_r134 = 32'b010001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane7_r134 = 32'b010001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane8_r134 = 32'b010001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane9_r134 = 32'b010001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane10_r134 = 32'b010001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane11_r134 = 32'b010001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane12_r134 = 32'b010001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane13_r134 = 32'b010001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane14_r134 = 32'b010001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane15_r134 = 32'b010001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane16_r134 = 32'b010001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane17_r134 = 32'b010001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane18_r134 = 32'b010001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane19_r134 = 32'b010001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane20_r134 = 32'b010001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane21_r134 = 32'b010001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane22_r134 = 32'b010001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane23_r134 = 32'b010001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane24_r134 = 32'b010001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane25_r134 = 32'b010001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane26_r134 = 32'b010001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane27_r134 = 32'b010001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane28_r134 = 32'b010001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane29_r134 = 32'b010001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane30_r134 = 32'b010001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.lane31_r134 = 32'b010001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[17].pe.lane0_r135 = 32'b010001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane1_r135 = 32'b010001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane2_r135 = 32'b010001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane3_r135 = 32'b010001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane4_r135 = 32'b010001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane5_r135 = 32'b010001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane6_r135 = 32'b010001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane7_r135 = 32'b010001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane8_r135 = 32'b010001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane9_r135 = 32'b010001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane10_r135 = 32'b010001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane11_r135 = 32'b010001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane12_r135 = 32'b010001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane13_r135 = 32'b010001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane14_r135 = 32'b010001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane15_r135 = 32'b010001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane16_r135 = 32'b010001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane17_r135 = 32'b010001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane18_r135 = 32'b010001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane19_r135 = 32'b010001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane20_r135 = 32'b010001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane21_r135 = 32'b010001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane22_r135 = 32'b010001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane23_r135 = 32'b010001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane24_r135 = 32'b010001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane25_r135 = 32'b010001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane26_r135 = 32'b010001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane27_r135 = 32'b010001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane28_r135 = 32'b010001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane29_r135 = 32'b010001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane30_r135 = 32'b010001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.lane31_r135 = 32'b010001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[18].pe.lane0_r134 = 32'b010010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane1_r134 = 32'b010010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane2_r134 = 32'b010010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane3_r134 = 32'b010010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane4_r134 = 32'b010010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane5_r134 = 32'b010010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane6_r134 = 32'b010010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane7_r134 = 32'b010010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane8_r134 = 32'b010010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane9_r134 = 32'b010010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane10_r134 = 32'b010010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane11_r134 = 32'b010010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane12_r134 = 32'b010010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane13_r134 = 32'b010010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane14_r134 = 32'b010010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane15_r134 = 32'b010010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane16_r134 = 32'b010010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane17_r134 = 32'b010010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane18_r134 = 32'b010010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane19_r134 = 32'b010010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane20_r134 = 32'b010010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane21_r134 = 32'b010010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane22_r134 = 32'b010010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane23_r134 = 32'b010010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane24_r134 = 32'b010010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane25_r134 = 32'b010010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane26_r134 = 32'b010010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane27_r134 = 32'b010010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane28_r134 = 32'b010010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane29_r134 = 32'b010010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane30_r134 = 32'b010010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.lane31_r134 = 32'b010010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[18].pe.lane0_r135 = 32'b010010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane1_r135 = 32'b010010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane2_r135 = 32'b010010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane3_r135 = 32'b010010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane4_r135 = 32'b010010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane5_r135 = 32'b010010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane6_r135 = 32'b010010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane7_r135 = 32'b010010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane8_r135 = 32'b010010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane9_r135 = 32'b010010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane10_r135 = 32'b010010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane11_r135 = 32'b010010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane12_r135 = 32'b010010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane13_r135 = 32'b010010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane14_r135 = 32'b010010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane15_r135 = 32'b010010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane16_r135 = 32'b010010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane17_r135 = 32'b010010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane18_r135 = 32'b010010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane19_r135 = 32'b010010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane20_r135 = 32'b010010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane21_r135 = 32'b010010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane22_r135 = 32'b010010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane23_r135 = 32'b010010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane24_r135 = 32'b010010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane25_r135 = 32'b010010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane26_r135 = 32'b010010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane27_r135 = 32'b010010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane28_r135 = 32'b010010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane29_r135 = 32'b010010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane30_r135 = 32'b010010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.lane31_r135 = 32'b010010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[19].pe.lane0_r134 = 32'b010011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane1_r134 = 32'b010011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane2_r134 = 32'b010011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane3_r134 = 32'b010011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane4_r134 = 32'b010011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane5_r134 = 32'b010011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane6_r134 = 32'b010011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane7_r134 = 32'b010011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane8_r134 = 32'b010011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane9_r134 = 32'b010011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane10_r134 = 32'b010011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane11_r134 = 32'b010011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane12_r134 = 32'b010011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane13_r134 = 32'b010011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane14_r134 = 32'b010011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane15_r134 = 32'b010011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane16_r134 = 32'b010011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane17_r134 = 32'b010011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane18_r134 = 32'b010011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane19_r134 = 32'b010011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane20_r134 = 32'b010011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane21_r134 = 32'b010011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane22_r134 = 32'b010011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane23_r134 = 32'b010011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane24_r134 = 32'b010011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane25_r134 = 32'b010011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane26_r134 = 32'b010011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane27_r134 = 32'b010011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane28_r134 = 32'b010011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane29_r134 = 32'b010011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane30_r134 = 32'b010011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.lane31_r134 = 32'b010011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[19].pe.lane0_r135 = 32'b010011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane1_r135 = 32'b010011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane2_r135 = 32'b010011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane3_r135 = 32'b010011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane4_r135 = 32'b010011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane5_r135 = 32'b010011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane6_r135 = 32'b010011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane7_r135 = 32'b010011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane8_r135 = 32'b010011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane9_r135 = 32'b010011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane10_r135 = 32'b010011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane11_r135 = 32'b010011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane12_r135 = 32'b010011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane13_r135 = 32'b010011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane14_r135 = 32'b010011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane15_r135 = 32'b010011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane16_r135 = 32'b010011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane17_r135 = 32'b010011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane18_r135 = 32'b010011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane19_r135 = 32'b010011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane20_r135 = 32'b010011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane21_r135 = 32'b010011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane22_r135 = 32'b010011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane23_r135 = 32'b010011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane24_r135 = 32'b010011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane25_r135 = 32'b010011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane26_r135 = 32'b010011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane27_r135 = 32'b010011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane28_r135 = 32'b010011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane29_r135 = 32'b010011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane30_r135 = 32'b010011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.lane31_r135 = 32'b010011_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[20].pe.lane0_r134 = 32'b010100_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane1_r134 = 32'b010100_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane2_r134 = 32'b010100_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane3_r134 = 32'b010100_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane4_r134 = 32'b010100_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane5_r134 = 32'b010100_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane6_r134 = 32'b010100_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane7_r134 = 32'b010100_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane8_r134 = 32'b010100_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane9_r134 = 32'b010100_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane10_r134 = 32'b010100_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane11_r134 = 32'b010100_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane12_r134 = 32'b010100_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane13_r134 = 32'b010100_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane14_r134 = 32'b010100_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane15_r134 = 32'b010100_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane16_r134 = 32'b010100_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane17_r134 = 32'b010100_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane18_r134 = 32'b010100_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane19_r134 = 32'b010100_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane20_r134 = 32'b010100_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane21_r134 = 32'b010100_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane22_r134 = 32'b010100_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane23_r134 = 32'b010100_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane24_r134 = 32'b010100_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane25_r134 = 32'b010100_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane26_r134 = 32'b010100_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane27_r134 = 32'b010100_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane28_r134 = 32'b010100_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane29_r134 = 32'b010100_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane30_r134 = 32'b010100_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.lane31_r134 = 32'b010100_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[20].pe.lane0_r135 = 32'b010100_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane1_r135 = 32'b010100_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane2_r135 = 32'b010100_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane3_r135 = 32'b010100_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane4_r135 = 32'b010100_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane5_r135 = 32'b010100_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane6_r135 = 32'b010100_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane7_r135 = 32'b010100_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane8_r135 = 32'b010100_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane9_r135 = 32'b010100_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane10_r135 = 32'b010100_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane11_r135 = 32'b010100_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane12_r135 = 32'b010100_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane13_r135 = 32'b010100_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane14_r135 = 32'b010100_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane15_r135 = 32'b010100_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane16_r135 = 32'b010100_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane17_r135 = 32'b010100_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane18_r135 = 32'b010100_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane19_r135 = 32'b010100_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane20_r135 = 32'b010100_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane21_r135 = 32'b010100_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane22_r135 = 32'b010100_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane23_r135 = 32'b010100_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane24_r135 = 32'b010100_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane25_r135 = 32'b010100_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane26_r135 = 32'b010100_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane27_r135 = 32'b010100_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane28_r135 = 32'b010100_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane29_r135 = 32'b010100_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane30_r135 = 32'b010100_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.lane31_r135 = 32'b010100_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[21].pe.lane0_r134 = 32'b010101_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane1_r134 = 32'b010101_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane2_r134 = 32'b010101_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane3_r134 = 32'b010101_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane4_r134 = 32'b010101_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane5_r134 = 32'b010101_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane6_r134 = 32'b010101_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane7_r134 = 32'b010101_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane8_r134 = 32'b010101_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane9_r134 = 32'b010101_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane10_r134 = 32'b010101_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane11_r134 = 32'b010101_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane12_r134 = 32'b010101_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane13_r134 = 32'b010101_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane14_r134 = 32'b010101_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane15_r134 = 32'b010101_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane16_r134 = 32'b010101_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane17_r134 = 32'b010101_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane18_r134 = 32'b010101_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane19_r134 = 32'b010101_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane20_r134 = 32'b010101_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane21_r134 = 32'b010101_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane22_r134 = 32'b010101_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane23_r134 = 32'b010101_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane24_r134 = 32'b010101_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane25_r134 = 32'b010101_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane26_r134 = 32'b010101_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane27_r134 = 32'b010101_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane28_r134 = 32'b010101_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane29_r134 = 32'b010101_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane30_r134 = 32'b010101_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.lane31_r134 = 32'b010101_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[21].pe.lane0_r135 = 32'b010101_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane1_r135 = 32'b010101_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane2_r135 = 32'b010101_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane3_r135 = 32'b010101_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane4_r135 = 32'b010101_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane5_r135 = 32'b010101_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane6_r135 = 32'b010101_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane7_r135 = 32'b010101_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane8_r135 = 32'b010101_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane9_r135 = 32'b010101_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane10_r135 = 32'b010101_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane11_r135 = 32'b010101_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane12_r135 = 32'b010101_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane13_r135 = 32'b010101_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane14_r135 = 32'b010101_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane15_r135 = 32'b010101_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane16_r135 = 32'b010101_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane17_r135 = 32'b010101_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane18_r135 = 32'b010101_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane19_r135 = 32'b010101_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane20_r135 = 32'b010101_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane21_r135 = 32'b010101_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane22_r135 = 32'b010101_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane23_r135 = 32'b010101_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane24_r135 = 32'b010101_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane25_r135 = 32'b010101_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane26_r135 = 32'b010101_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane27_r135 = 32'b010101_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane28_r135 = 32'b010101_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane29_r135 = 32'b010101_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane30_r135 = 32'b010101_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.lane31_r135 = 32'b010101_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[22].pe.lane0_r134 = 32'b010110_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane1_r134 = 32'b010110_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane2_r134 = 32'b010110_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane3_r134 = 32'b010110_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane4_r134 = 32'b010110_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane5_r134 = 32'b010110_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane6_r134 = 32'b010110_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane7_r134 = 32'b010110_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane8_r134 = 32'b010110_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane9_r134 = 32'b010110_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane10_r134 = 32'b010110_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane11_r134 = 32'b010110_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane12_r134 = 32'b010110_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane13_r134 = 32'b010110_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane14_r134 = 32'b010110_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane15_r134 = 32'b010110_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane16_r134 = 32'b010110_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane17_r134 = 32'b010110_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane18_r134 = 32'b010110_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane19_r134 = 32'b010110_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane20_r134 = 32'b010110_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane21_r134 = 32'b010110_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane22_r134 = 32'b010110_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane23_r134 = 32'b010110_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane24_r134 = 32'b010110_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane25_r134 = 32'b010110_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane26_r134 = 32'b010110_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane27_r134 = 32'b010110_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane28_r134 = 32'b010110_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane29_r134 = 32'b010110_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane30_r134 = 32'b010110_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.lane31_r134 = 32'b010110_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[22].pe.lane0_r135 = 32'b010110_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane1_r135 = 32'b010110_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane2_r135 = 32'b010110_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane3_r135 = 32'b010110_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane4_r135 = 32'b010110_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane5_r135 = 32'b010110_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane6_r135 = 32'b010110_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane7_r135 = 32'b010110_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane8_r135 = 32'b010110_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane9_r135 = 32'b010110_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane10_r135 = 32'b010110_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane11_r135 = 32'b010110_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane12_r135 = 32'b010110_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane13_r135 = 32'b010110_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane14_r135 = 32'b010110_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane15_r135 = 32'b010110_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane16_r135 = 32'b010110_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane17_r135 = 32'b010110_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane18_r135 = 32'b010110_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane19_r135 = 32'b010110_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane20_r135 = 32'b010110_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane21_r135 = 32'b010110_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane22_r135 = 32'b010110_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane23_r135 = 32'b010110_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane24_r135 = 32'b010110_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane25_r135 = 32'b010110_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane26_r135 = 32'b010110_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane27_r135 = 32'b010110_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane28_r135 = 32'b010110_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane29_r135 = 32'b010110_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane30_r135 = 32'b010110_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.lane31_r135 = 32'b010110_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[23].pe.lane0_r134 = 32'b010111_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane1_r134 = 32'b010111_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane2_r134 = 32'b010111_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane3_r134 = 32'b010111_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane4_r134 = 32'b010111_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane5_r134 = 32'b010111_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane6_r134 = 32'b010111_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane7_r134 = 32'b010111_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane8_r134 = 32'b010111_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane9_r134 = 32'b010111_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane10_r134 = 32'b010111_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane11_r134 = 32'b010111_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane12_r134 = 32'b010111_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane13_r134 = 32'b010111_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane14_r134 = 32'b010111_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane15_r134 = 32'b010111_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane16_r134 = 32'b010111_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane17_r134 = 32'b010111_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane18_r134 = 32'b010111_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane19_r134 = 32'b010111_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane20_r134 = 32'b010111_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane21_r134 = 32'b010111_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane22_r134 = 32'b010111_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane23_r134 = 32'b010111_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane24_r134 = 32'b010111_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane25_r134 = 32'b010111_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane26_r134 = 32'b010111_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane27_r134 = 32'b010111_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane28_r134 = 32'b010111_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane29_r134 = 32'b010111_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane30_r134 = 32'b010111_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.lane31_r134 = 32'b010111_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[23].pe.lane0_r135 = 32'b010111_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane1_r135 = 32'b010111_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane2_r135 = 32'b010111_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane3_r135 = 32'b010111_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane4_r135 = 32'b010111_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane5_r135 = 32'b010111_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane6_r135 = 32'b010111_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane7_r135 = 32'b010111_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane8_r135 = 32'b010111_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane9_r135 = 32'b010111_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane10_r135 = 32'b010111_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane11_r135 = 32'b010111_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane12_r135 = 32'b010111_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane13_r135 = 32'b010111_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane14_r135 = 32'b010111_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane15_r135 = 32'b010111_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane16_r135 = 32'b010111_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane17_r135 = 32'b010111_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane18_r135 = 32'b010111_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane19_r135 = 32'b010111_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane20_r135 = 32'b010111_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane21_r135 = 32'b010111_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane22_r135 = 32'b010111_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane23_r135 = 32'b010111_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane24_r135 = 32'b010111_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane25_r135 = 32'b010111_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane26_r135 = 32'b010111_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane27_r135 = 32'b010111_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane28_r135 = 32'b010111_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane29_r135 = 32'b010111_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane30_r135 = 32'b010111_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.lane31_r135 = 32'b010111_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[24].pe.lane0_r134 = 32'b011000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane1_r134 = 32'b011000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane2_r134 = 32'b011000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane3_r134 = 32'b011000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane4_r134 = 32'b011000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane5_r134 = 32'b011000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane6_r134 = 32'b011000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane7_r134 = 32'b011000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane8_r134 = 32'b011000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane9_r134 = 32'b011000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane10_r134 = 32'b011000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane11_r134 = 32'b011000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane12_r134 = 32'b011000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane13_r134 = 32'b011000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane14_r134 = 32'b011000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane15_r134 = 32'b011000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane16_r134 = 32'b011000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane17_r134 = 32'b011000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane18_r134 = 32'b011000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane19_r134 = 32'b011000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane20_r134 = 32'b011000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane21_r134 = 32'b011000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane22_r134 = 32'b011000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane23_r134 = 32'b011000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane24_r134 = 32'b011000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane25_r134 = 32'b011000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane26_r134 = 32'b011000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane27_r134 = 32'b011000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane28_r134 = 32'b011000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane29_r134 = 32'b011000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane30_r134 = 32'b011000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.lane31_r134 = 32'b011000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[24].pe.lane0_r135 = 32'b011000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane1_r135 = 32'b011000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane2_r135 = 32'b011000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane3_r135 = 32'b011000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane4_r135 = 32'b011000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane5_r135 = 32'b011000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane6_r135 = 32'b011000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane7_r135 = 32'b011000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane8_r135 = 32'b011000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane9_r135 = 32'b011000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane10_r135 = 32'b011000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane11_r135 = 32'b011000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane12_r135 = 32'b011000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane13_r135 = 32'b011000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane14_r135 = 32'b011000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane15_r135 = 32'b011000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane16_r135 = 32'b011000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane17_r135 = 32'b011000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane18_r135 = 32'b011000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane19_r135 = 32'b011000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane20_r135 = 32'b011000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane21_r135 = 32'b011000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane22_r135 = 32'b011000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane23_r135 = 32'b011000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane24_r135 = 32'b011000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane25_r135 = 32'b011000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane26_r135 = 32'b011000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane27_r135 = 32'b011000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane28_r135 = 32'b011000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane29_r135 = 32'b011000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane30_r135 = 32'b011000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.lane31_r135 = 32'b011000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[25].pe.lane0_r134 = 32'b011001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane1_r134 = 32'b011001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane2_r134 = 32'b011001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane3_r134 = 32'b011001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane4_r134 = 32'b011001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane5_r134 = 32'b011001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane6_r134 = 32'b011001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane7_r134 = 32'b011001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane8_r134 = 32'b011001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane9_r134 = 32'b011001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane10_r134 = 32'b011001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane11_r134 = 32'b011001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane12_r134 = 32'b011001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane13_r134 = 32'b011001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane14_r134 = 32'b011001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane15_r134 = 32'b011001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane16_r134 = 32'b011001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane17_r134 = 32'b011001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane18_r134 = 32'b011001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane19_r134 = 32'b011001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane20_r134 = 32'b011001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane21_r134 = 32'b011001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane22_r134 = 32'b011001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane23_r134 = 32'b011001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane24_r134 = 32'b011001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane25_r134 = 32'b011001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane26_r134 = 32'b011001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane27_r134 = 32'b011001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane28_r134 = 32'b011001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane29_r134 = 32'b011001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane30_r134 = 32'b011001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.lane31_r134 = 32'b011001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[25].pe.lane0_r135 = 32'b011001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane1_r135 = 32'b011001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane2_r135 = 32'b011001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane3_r135 = 32'b011001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane4_r135 = 32'b011001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane5_r135 = 32'b011001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane6_r135 = 32'b011001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane7_r135 = 32'b011001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane8_r135 = 32'b011001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane9_r135 = 32'b011001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane10_r135 = 32'b011001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane11_r135 = 32'b011001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane12_r135 = 32'b011001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane13_r135 = 32'b011001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane14_r135 = 32'b011001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane15_r135 = 32'b011001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane16_r135 = 32'b011001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane17_r135 = 32'b011001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane18_r135 = 32'b011001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane19_r135 = 32'b011001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane20_r135 = 32'b011001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane21_r135 = 32'b011001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane22_r135 = 32'b011001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane23_r135 = 32'b011001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane24_r135 = 32'b011001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane25_r135 = 32'b011001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane26_r135 = 32'b011001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane27_r135 = 32'b011001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane28_r135 = 32'b011001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane29_r135 = 32'b011001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane30_r135 = 32'b011001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.lane31_r135 = 32'b011001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[26].pe.lane0_r134 = 32'b011010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane1_r134 = 32'b011010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane2_r134 = 32'b011010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane3_r134 = 32'b011010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane4_r134 = 32'b011010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane5_r134 = 32'b011010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane6_r134 = 32'b011010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane7_r134 = 32'b011010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane8_r134 = 32'b011010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane9_r134 = 32'b011010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane10_r134 = 32'b011010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane11_r134 = 32'b011010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane12_r134 = 32'b011010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane13_r134 = 32'b011010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane14_r134 = 32'b011010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane15_r134 = 32'b011010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane16_r134 = 32'b011010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane17_r134 = 32'b011010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane18_r134 = 32'b011010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane19_r134 = 32'b011010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane20_r134 = 32'b011010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane21_r134 = 32'b011010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane22_r134 = 32'b011010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane23_r134 = 32'b011010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane24_r134 = 32'b011010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane25_r134 = 32'b011010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane26_r134 = 32'b011010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane27_r134 = 32'b011010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane28_r134 = 32'b011010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane29_r134 = 32'b011010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane30_r134 = 32'b011010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.lane31_r134 = 32'b011010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[26].pe.lane0_r135 = 32'b011010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane1_r135 = 32'b011010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane2_r135 = 32'b011010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane3_r135 = 32'b011010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane4_r135 = 32'b011010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane5_r135 = 32'b011010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane6_r135 = 32'b011010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane7_r135 = 32'b011010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane8_r135 = 32'b011010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane9_r135 = 32'b011010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane10_r135 = 32'b011010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane11_r135 = 32'b011010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane12_r135 = 32'b011010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane13_r135 = 32'b011010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane14_r135 = 32'b011010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane15_r135 = 32'b011010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane16_r135 = 32'b011010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane17_r135 = 32'b011010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane18_r135 = 32'b011010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane19_r135 = 32'b011010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane20_r135 = 32'b011010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane21_r135 = 32'b011010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane22_r135 = 32'b011010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane23_r135 = 32'b011010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane24_r135 = 32'b011010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane25_r135 = 32'b011010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane26_r135 = 32'b011010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane27_r135 = 32'b011010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane28_r135 = 32'b011010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane29_r135 = 32'b011010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane30_r135 = 32'b011010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.lane31_r135 = 32'b011010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[27].pe.lane0_r134 = 32'b011011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane1_r134 = 32'b011011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane2_r134 = 32'b011011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane3_r134 = 32'b011011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane4_r134 = 32'b011011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane5_r134 = 32'b011011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane6_r134 = 32'b011011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane7_r134 = 32'b011011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane8_r134 = 32'b011011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane9_r134 = 32'b011011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane10_r134 = 32'b011011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane11_r134 = 32'b011011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane12_r134 = 32'b011011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane13_r134 = 32'b011011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane14_r134 = 32'b011011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane15_r134 = 32'b011011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane16_r134 = 32'b011011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane17_r134 = 32'b011011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane18_r134 = 32'b011011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane19_r134 = 32'b011011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane20_r134 = 32'b011011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane21_r134 = 32'b011011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane22_r134 = 32'b011011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane23_r134 = 32'b011011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane24_r134 = 32'b011011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane25_r134 = 32'b011011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane26_r134 = 32'b011011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane27_r134 = 32'b011011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane28_r134 = 32'b011011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane29_r134 = 32'b011011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane30_r134 = 32'b011011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.lane31_r134 = 32'b011011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[27].pe.lane0_r135 = 32'b011011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane1_r135 = 32'b011011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane2_r135 = 32'b011011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane3_r135 = 32'b011011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane4_r135 = 32'b011011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane5_r135 = 32'b011011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane6_r135 = 32'b011011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane7_r135 = 32'b011011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane8_r135 = 32'b011011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane9_r135 = 32'b011011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane10_r135 = 32'b011011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane11_r135 = 32'b011011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane12_r135 = 32'b011011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane13_r135 = 32'b011011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane14_r135 = 32'b011011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane15_r135 = 32'b011011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane16_r135 = 32'b011011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane17_r135 = 32'b011011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane18_r135 = 32'b011011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane19_r135 = 32'b011011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane20_r135 = 32'b011011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane21_r135 = 32'b011011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane22_r135 = 32'b011011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane23_r135 = 32'b011011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane24_r135 = 32'b011011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane25_r135 = 32'b011011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane26_r135 = 32'b011011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane27_r135 = 32'b011011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane28_r135 = 32'b011011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane29_r135 = 32'b011011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane30_r135 = 32'b011011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.lane31_r135 = 32'b011011_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[28].pe.lane0_r134 = 32'b011100_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane1_r134 = 32'b011100_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane2_r134 = 32'b011100_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane3_r134 = 32'b011100_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane4_r134 = 32'b011100_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane5_r134 = 32'b011100_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane6_r134 = 32'b011100_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane7_r134 = 32'b011100_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane8_r134 = 32'b011100_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane9_r134 = 32'b011100_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane10_r134 = 32'b011100_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane11_r134 = 32'b011100_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane12_r134 = 32'b011100_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane13_r134 = 32'b011100_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane14_r134 = 32'b011100_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane15_r134 = 32'b011100_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane16_r134 = 32'b011100_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane17_r134 = 32'b011100_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane18_r134 = 32'b011100_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane19_r134 = 32'b011100_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane20_r134 = 32'b011100_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane21_r134 = 32'b011100_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane22_r134 = 32'b011100_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane23_r134 = 32'b011100_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane24_r134 = 32'b011100_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane25_r134 = 32'b011100_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane26_r134 = 32'b011100_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane27_r134 = 32'b011100_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane28_r134 = 32'b011100_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane29_r134 = 32'b011100_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane30_r134 = 32'b011100_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.lane31_r134 = 32'b011100_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[28].pe.lane0_r135 = 32'b011100_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane1_r135 = 32'b011100_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane2_r135 = 32'b011100_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane3_r135 = 32'b011100_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane4_r135 = 32'b011100_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane5_r135 = 32'b011100_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane6_r135 = 32'b011100_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane7_r135 = 32'b011100_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane8_r135 = 32'b011100_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane9_r135 = 32'b011100_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane10_r135 = 32'b011100_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane11_r135 = 32'b011100_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane12_r135 = 32'b011100_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane13_r135 = 32'b011100_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane14_r135 = 32'b011100_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane15_r135 = 32'b011100_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane16_r135 = 32'b011100_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane17_r135 = 32'b011100_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane18_r135 = 32'b011100_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane19_r135 = 32'b011100_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane20_r135 = 32'b011100_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane21_r135 = 32'b011100_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane22_r135 = 32'b011100_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane23_r135 = 32'b011100_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane24_r135 = 32'b011100_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane25_r135 = 32'b011100_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane26_r135 = 32'b011100_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane27_r135 = 32'b011100_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane28_r135 = 32'b011100_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane29_r135 = 32'b011100_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane30_r135 = 32'b011100_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.lane31_r135 = 32'b011100_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[29].pe.lane0_r134 = 32'b011101_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane1_r134 = 32'b011101_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane2_r134 = 32'b011101_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane3_r134 = 32'b011101_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane4_r134 = 32'b011101_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane5_r134 = 32'b011101_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane6_r134 = 32'b011101_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane7_r134 = 32'b011101_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane8_r134 = 32'b011101_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane9_r134 = 32'b011101_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane10_r134 = 32'b011101_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane11_r134 = 32'b011101_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane12_r134 = 32'b011101_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane13_r134 = 32'b011101_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane14_r134 = 32'b011101_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane15_r134 = 32'b011101_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane16_r134 = 32'b011101_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane17_r134 = 32'b011101_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane18_r134 = 32'b011101_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane19_r134 = 32'b011101_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane20_r134 = 32'b011101_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane21_r134 = 32'b011101_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane22_r134 = 32'b011101_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane23_r134 = 32'b011101_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane24_r134 = 32'b011101_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane25_r134 = 32'b011101_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane26_r134 = 32'b011101_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane27_r134 = 32'b011101_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane28_r134 = 32'b011101_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane29_r134 = 32'b011101_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane30_r134 = 32'b011101_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.lane31_r134 = 32'b011101_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[29].pe.lane0_r135 = 32'b011101_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane1_r135 = 32'b011101_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane2_r135 = 32'b011101_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane3_r135 = 32'b011101_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane4_r135 = 32'b011101_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane5_r135 = 32'b011101_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane6_r135 = 32'b011101_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane7_r135 = 32'b011101_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane8_r135 = 32'b011101_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane9_r135 = 32'b011101_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane10_r135 = 32'b011101_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane11_r135 = 32'b011101_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane12_r135 = 32'b011101_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane13_r135 = 32'b011101_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane14_r135 = 32'b011101_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane15_r135 = 32'b011101_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane16_r135 = 32'b011101_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane17_r135 = 32'b011101_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane18_r135 = 32'b011101_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane19_r135 = 32'b011101_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane20_r135 = 32'b011101_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane21_r135 = 32'b011101_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane22_r135 = 32'b011101_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane23_r135 = 32'b011101_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane24_r135 = 32'b011101_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane25_r135 = 32'b011101_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane26_r135 = 32'b011101_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane27_r135 = 32'b011101_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane28_r135 = 32'b011101_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane29_r135 = 32'b011101_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane30_r135 = 32'b011101_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.lane31_r135 = 32'b011101_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[30].pe.lane0_r134 = 32'b011110_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane1_r134 = 32'b011110_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane2_r134 = 32'b011110_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane3_r134 = 32'b011110_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane4_r134 = 32'b011110_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane5_r134 = 32'b011110_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane6_r134 = 32'b011110_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane7_r134 = 32'b011110_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane8_r134 = 32'b011110_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane9_r134 = 32'b011110_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane10_r134 = 32'b011110_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane11_r134 = 32'b011110_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane12_r134 = 32'b011110_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane13_r134 = 32'b011110_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane14_r134 = 32'b011110_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane15_r134 = 32'b011110_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane16_r134 = 32'b011110_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane17_r134 = 32'b011110_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane18_r134 = 32'b011110_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane19_r134 = 32'b011110_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane20_r134 = 32'b011110_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane21_r134 = 32'b011110_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane22_r134 = 32'b011110_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane23_r134 = 32'b011110_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane24_r134 = 32'b011110_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane25_r134 = 32'b011110_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane26_r134 = 32'b011110_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane27_r134 = 32'b011110_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane28_r134 = 32'b011110_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane29_r134 = 32'b011110_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane30_r134 = 32'b011110_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.lane31_r134 = 32'b011110_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[30].pe.lane0_r135 = 32'b011110_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane1_r135 = 32'b011110_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane2_r135 = 32'b011110_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane3_r135 = 32'b011110_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane4_r135 = 32'b011110_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane5_r135 = 32'b011110_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane6_r135 = 32'b011110_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane7_r135 = 32'b011110_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane8_r135 = 32'b011110_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane9_r135 = 32'b011110_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane10_r135 = 32'b011110_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane11_r135 = 32'b011110_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane12_r135 = 32'b011110_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane13_r135 = 32'b011110_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane14_r135 = 32'b011110_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane15_r135 = 32'b011110_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane16_r135 = 32'b011110_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane17_r135 = 32'b011110_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane18_r135 = 32'b011110_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane19_r135 = 32'b011110_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane20_r135 = 32'b011110_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane21_r135 = 32'b011110_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane22_r135 = 32'b011110_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane23_r135 = 32'b011110_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane24_r135 = 32'b011110_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane25_r135 = 32'b011110_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane26_r135 = 32'b011110_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane27_r135 = 32'b011110_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane28_r135 = 32'b011110_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane29_r135 = 32'b011110_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane30_r135 = 32'b011110_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.lane31_r135 = 32'b011110_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[31].pe.lane0_r134 = 32'b011111_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane1_r134 = 32'b011111_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane2_r134 = 32'b011111_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane3_r134 = 32'b011111_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane4_r134 = 32'b011111_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane5_r134 = 32'b011111_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane6_r134 = 32'b011111_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane7_r134 = 32'b011111_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane8_r134 = 32'b011111_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane9_r134 = 32'b011111_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane10_r134 = 32'b011111_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane11_r134 = 32'b011111_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane12_r134 = 32'b011111_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane13_r134 = 32'b011111_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane14_r134 = 32'b011111_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane15_r134 = 32'b011111_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane16_r134 = 32'b011111_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane17_r134 = 32'b011111_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane18_r134 = 32'b011111_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane19_r134 = 32'b011111_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane20_r134 = 32'b011111_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane21_r134 = 32'b011111_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane22_r134 = 32'b011111_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane23_r134 = 32'b011111_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane24_r134 = 32'b011111_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane25_r134 = 32'b011111_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane26_r134 = 32'b011111_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane27_r134 = 32'b011111_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane28_r134 = 32'b011111_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane29_r134 = 32'b011111_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane30_r134 = 32'b011111_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.lane31_r134 = 32'b011111_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[31].pe.lane0_r135 = 32'b011111_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane1_r135 = 32'b011111_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane2_r135 = 32'b011111_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane3_r135 = 32'b011111_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane4_r135 = 32'b011111_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane5_r135 = 32'b011111_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane6_r135 = 32'b011111_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane7_r135 = 32'b011111_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane8_r135 = 32'b011111_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane9_r135 = 32'b011111_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane10_r135 = 32'b011111_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane11_r135 = 32'b011111_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane12_r135 = 32'b011111_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane13_r135 = 32'b011111_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane14_r135 = 32'b011111_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane15_r135 = 32'b011111_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane16_r135 = 32'b011111_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane17_r135 = 32'b011111_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane18_r135 = 32'b011111_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane19_r135 = 32'b011111_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane20_r135 = 32'b011111_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane21_r135 = 32'b011111_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane22_r135 = 32'b011111_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane23_r135 = 32'b011111_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane24_r135 = 32'b011111_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane25_r135 = 32'b011111_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane26_r135 = 32'b011111_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane27_r135 = 32'b011111_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane28_r135 = 32'b011111_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane29_r135 = 32'b011111_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane30_r135 = 32'b011111_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.lane31_r135 = 32'b011111_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[32].pe.lane0_r134 = 32'b100000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane1_r134 = 32'b100000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane2_r134 = 32'b100000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane3_r134 = 32'b100000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane4_r134 = 32'b100000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane5_r134 = 32'b100000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane6_r134 = 32'b100000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane7_r134 = 32'b100000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane8_r134 = 32'b100000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane9_r134 = 32'b100000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane10_r134 = 32'b100000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane11_r134 = 32'b100000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane12_r134 = 32'b100000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane13_r134 = 32'b100000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane14_r134 = 32'b100000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane15_r134 = 32'b100000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane16_r134 = 32'b100000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane17_r134 = 32'b100000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane18_r134 = 32'b100000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane19_r134 = 32'b100000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane20_r134 = 32'b100000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane21_r134 = 32'b100000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane22_r134 = 32'b100000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane23_r134 = 32'b100000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane24_r134 = 32'b100000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane25_r134 = 32'b100000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane26_r134 = 32'b100000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane27_r134 = 32'b100000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane28_r134 = 32'b100000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane29_r134 = 32'b100000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane30_r134 = 32'b100000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.lane31_r134 = 32'b100000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[32].pe.lane0_r135 = 32'b100000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane1_r135 = 32'b100000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane2_r135 = 32'b100000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane3_r135 = 32'b100000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane4_r135 = 32'b100000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane5_r135 = 32'b100000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane6_r135 = 32'b100000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane7_r135 = 32'b100000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane8_r135 = 32'b100000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane9_r135 = 32'b100000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane10_r135 = 32'b100000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane11_r135 = 32'b100000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane12_r135 = 32'b100000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane13_r135 = 32'b100000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane14_r135 = 32'b100000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane15_r135 = 32'b100000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane16_r135 = 32'b100000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane17_r135 = 32'b100000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane18_r135 = 32'b100000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane19_r135 = 32'b100000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane20_r135 = 32'b100000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane21_r135 = 32'b100000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane22_r135 = 32'b100000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane23_r135 = 32'b100000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane24_r135 = 32'b100000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane25_r135 = 32'b100000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane26_r135 = 32'b100000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane27_r135 = 32'b100000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane28_r135 = 32'b100000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane29_r135 = 32'b100000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane30_r135 = 32'b100000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.lane31_r135 = 32'b100000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[33].pe.lane0_r134 = 32'b100001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane1_r134 = 32'b100001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane2_r134 = 32'b100001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane3_r134 = 32'b100001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane4_r134 = 32'b100001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane5_r134 = 32'b100001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane6_r134 = 32'b100001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane7_r134 = 32'b100001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane8_r134 = 32'b100001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane9_r134 = 32'b100001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane10_r134 = 32'b100001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane11_r134 = 32'b100001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane12_r134 = 32'b100001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane13_r134 = 32'b100001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane14_r134 = 32'b100001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane15_r134 = 32'b100001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane16_r134 = 32'b100001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane17_r134 = 32'b100001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane18_r134 = 32'b100001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane19_r134 = 32'b100001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane20_r134 = 32'b100001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane21_r134 = 32'b100001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane22_r134 = 32'b100001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane23_r134 = 32'b100001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane24_r134 = 32'b100001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane25_r134 = 32'b100001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane26_r134 = 32'b100001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane27_r134 = 32'b100001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane28_r134 = 32'b100001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane29_r134 = 32'b100001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane30_r134 = 32'b100001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.lane31_r134 = 32'b100001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[33].pe.lane0_r135 = 32'b100001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane1_r135 = 32'b100001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane2_r135 = 32'b100001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane3_r135 = 32'b100001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane4_r135 = 32'b100001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane5_r135 = 32'b100001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane6_r135 = 32'b100001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane7_r135 = 32'b100001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane8_r135 = 32'b100001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane9_r135 = 32'b100001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane10_r135 = 32'b100001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane11_r135 = 32'b100001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane12_r135 = 32'b100001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane13_r135 = 32'b100001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane14_r135 = 32'b100001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane15_r135 = 32'b100001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane16_r135 = 32'b100001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane17_r135 = 32'b100001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane18_r135 = 32'b100001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane19_r135 = 32'b100001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane20_r135 = 32'b100001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane21_r135 = 32'b100001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane22_r135 = 32'b100001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane23_r135 = 32'b100001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane24_r135 = 32'b100001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane25_r135 = 32'b100001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane26_r135 = 32'b100001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane27_r135 = 32'b100001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane28_r135 = 32'b100001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane29_r135 = 32'b100001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane30_r135 = 32'b100001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.lane31_r135 = 32'b100001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[34].pe.lane0_r134 = 32'b100010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane1_r134 = 32'b100010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane2_r134 = 32'b100010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane3_r134 = 32'b100010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane4_r134 = 32'b100010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane5_r134 = 32'b100010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane6_r134 = 32'b100010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane7_r134 = 32'b100010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane8_r134 = 32'b100010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane9_r134 = 32'b100010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane10_r134 = 32'b100010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane11_r134 = 32'b100010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane12_r134 = 32'b100010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane13_r134 = 32'b100010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane14_r134 = 32'b100010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane15_r134 = 32'b100010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane16_r134 = 32'b100010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane17_r134 = 32'b100010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane18_r134 = 32'b100010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane19_r134 = 32'b100010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane20_r134 = 32'b100010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane21_r134 = 32'b100010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane22_r134 = 32'b100010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane23_r134 = 32'b100010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane24_r134 = 32'b100010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane25_r134 = 32'b100010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane26_r134 = 32'b100010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane27_r134 = 32'b100010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane28_r134 = 32'b100010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane29_r134 = 32'b100010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane30_r134 = 32'b100010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.lane31_r134 = 32'b100010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[34].pe.lane0_r135 = 32'b100010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane1_r135 = 32'b100010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane2_r135 = 32'b100010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane3_r135 = 32'b100010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane4_r135 = 32'b100010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane5_r135 = 32'b100010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane6_r135 = 32'b100010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane7_r135 = 32'b100010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane8_r135 = 32'b100010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane9_r135 = 32'b100010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane10_r135 = 32'b100010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane11_r135 = 32'b100010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane12_r135 = 32'b100010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane13_r135 = 32'b100010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane14_r135 = 32'b100010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane15_r135 = 32'b100010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane16_r135 = 32'b100010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane17_r135 = 32'b100010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane18_r135 = 32'b100010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane19_r135 = 32'b100010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane20_r135 = 32'b100010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane21_r135 = 32'b100010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane22_r135 = 32'b100010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane23_r135 = 32'b100010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane24_r135 = 32'b100010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane25_r135 = 32'b100010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane26_r135 = 32'b100010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane27_r135 = 32'b100010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane28_r135 = 32'b100010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane29_r135 = 32'b100010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane30_r135 = 32'b100010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.lane31_r135 = 32'b100010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[35].pe.lane0_r134 = 32'b100011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane1_r134 = 32'b100011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane2_r134 = 32'b100011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane3_r134 = 32'b100011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane4_r134 = 32'b100011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane5_r134 = 32'b100011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane6_r134 = 32'b100011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane7_r134 = 32'b100011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane8_r134 = 32'b100011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane9_r134 = 32'b100011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane10_r134 = 32'b100011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane11_r134 = 32'b100011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane12_r134 = 32'b100011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane13_r134 = 32'b100011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane14_r134 = 32'b100011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane15_r134 = 32'b100011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane16_r134 = 32'b100011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane17_r134 = 32'b100011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane18_r134 = 32'b100011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane19_r134 = 32'b100011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane20_r134 = 32'b100011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane21_r134 = 32'b100011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane22_r134 = 32'b100011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane23_r134 = 32'b100011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane24_r134 = 32'b100011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane25_r134 = 32'b100011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane26_r134 = 32'b100011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane27_r134 = 32'b100011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane28_r134 = 32'b100011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane29_r134 = 32'b100011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane30_r134 = 32'b100011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.lane31_r134 = 32'b100011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[35].pe.lane0_r135 = 32'b100011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane1_r135 = 32'b100011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane2_r135 = 32'b100011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane3_r135 = 32'b100011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane4_r135 = 32'b100011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane5_r135 = 32'b100011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane6_r135 = 32'b100011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane7_r135 = 32'b100011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane8_r135 = 32'b100011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane9_r135 = 32'b100011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane10_r135 = 32'b100011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane11_r135 = 32'b100011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane12_r135 = 32'b100011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane13_r135 = 32'b100011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane14_r135 = 32'b100011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane15_r135 = 32'b100011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane16_r135 = 32'b100011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane17_r135 = 32'b100011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane18_r135 = 32'b100011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane19_r135 = 32'b100011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane20_r135 = 32'b100011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane21_r135 = 32'b100011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane22_r135 = 32'b100011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane23_r135 = 32'b100011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane24_r135 = 32'b100011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane25_r135 = 32'b100011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane26_r135 = 32'b100011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane27_r135 = 32'b100011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane28_r135 = 32'b100011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane29_r135 = 32'b100011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane30_r135 = 32'b100011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.lane31_r135 = 32'b100011_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[36].pe.lane0_r134 = 32'b100100_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane1_r134 = 32'b100100_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane2_r134 = 32'b100100_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane3_r134 = 32'b100100_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane4_r134 = 32'b100100_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane5_r134 = 32'b100100_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane6_r134 = 32'b100100_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane7_r134 = 32'b100100_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane8_r134 = 32'b100100_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane9_r134 = 32'b100100_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane10_r134 = 32'b100100_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane11_r134 = 32'b100100_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane12_r134 = 32'b100100_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane13_r134 = 32'b100100_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane14_r134 = 32'b100100_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane15_r134 = 32'b100100_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane16_r134 = 32'b100100_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane17_r134 = 32'b100100_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane18_r134 = 32'b100100_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane19_r134 = 32'b100100_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane20_r134 = 32'b100100_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane21_r134 = 32'b100100_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane22_r134 = 32'b100100_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane23_r134 = 32'b100100_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane24_r134 = 32'b100100_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane25_r134 = 32'b100100_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane26_r134 = 32'b100100_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane27_r134 = 32'b100100_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane28_r134 = 32'b100100_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane29_r134 = 32'b100100_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane30_r134 = 32'b100100_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.lane31_r134 = 32'b100100_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[36].pe.lane0_r135 = 32'b100100_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane1_r135 = 32'b100100_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane2_r135 = 32'b100100_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane3_r135 = 32'b100100_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane4_r135 = 32'b100100_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane5_r135 = 32'b100100_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane6_r135 = 32'b100100_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane7_r135 = 32'b100100_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane8_r135 = 32'b100100_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane9_r135 = 32'b100100_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane10_r135 = 32'b100100_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane11_r135 = 32'b100100_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane12_r135 = 32'b100100_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane13_r135 = 32'b100100_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane14_r135 = 32'b100100_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane15_r135 = 32'b100100_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane16_r135 = 32'b100100_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane17_r135 = 32'b100100_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane18_r135 = 32'b100100_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane19_r135 = 32'b100100_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane20_r135 = 32'b100100_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane21_r135 = 32'b100100_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane22_r135 = 32'b100100_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane23_r135 = 32'b100100_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane24_r135 = 32'b100100_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane25_r135 = 32'b100100_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane26_r135 = 32'b100100_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane27_r135 = 32'b100100_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane28_r135 = 32'b100100_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane29_r135 = 32'b100100_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane30_r135 = 32'b100100_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.lane31_r135 = 32'b100100_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[37].pe.lane0_r134 = 32'b100101_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane1_r134 = 32'b100101_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane2_r134 = 32'b100101_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane3_r134 = 32'b100101_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane4_r134 = 32'b100101_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane5_r134 = 32'b100101_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane6_r134 = 32'b100101_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane7_r134 = 32'b100101_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane8_r134 = 32'b100101_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane9_r134 = 32'b100101_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane10_r134 = 32'b100101_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane11_r134 = 32'b100101_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane12_r134 = 32'b100101_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane13_r134 = 32'b100101_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane14_r134 = 32'b100101_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane15_r134 = 32'b100101_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane16_r134 = 32'b100101_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane17_r134 = 32'b100101_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane18_r134 = 32'b100101_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane19_r134 = 32'b100101_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane20_r134 = 32'b100101_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane21_r134 = 32'b100101_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane22_r134 = 32'b100101_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane23_r134 = 32'b100101_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane24_r134 = 32'b100101_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane25_r134 = 32'b100101_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane26_r134 = 32'b100101_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane27_r134 = 32'b100101_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane28_r134 = 32'b100101_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane29_r134 = 32'b100101_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane30_r134 = 32'b100101_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.lane31_r134 = 32'b100101_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[37].pe.lane0_r135 = 32'b100101_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane1_r135 = 32'b100101_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane2_r135 = 32'b100101_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane3_r135 = 32'b100101_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane4_r135 = 32'b100101_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane5_r135 = 32'b100101_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane6_r135 = 32'b100101_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane7_r135 = 32'b100101_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane8_r135 = 32'b100101_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane9_r135 = 32'b100101_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane10_r135 = 32'b100101_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane11_r135 = 32'b100101_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane12_r135 = 32'b100101_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane13_r135 = 32'b100101_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane14_r135 = 32'b100101_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane15_r135 = 32'b100101_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane16_r135 = 32'b100101_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane17_r135 = 32'b100101_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane18_r135 = 32'b100101_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane19_r135 = 32'b100101_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane20_r135 = 32'b100101_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane21_r135 = 32'b100101_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane22_r135 = 32'b100101_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane23_r135 = 32'b100101_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane24_r135 = 32'b100101_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane25_r135 = 32'b100101_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane26_r135 = 32'b100101_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane27_r135 = 32'b100101_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane28_r135 = 32'b100101_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane29_r135 = 32'b100101_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane30_r135 = 32'b100101_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.lane31_r135 = 32'b100101_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[38].pe.lane0_r134 = 32'b100110_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane1_r134 = 32'b100110_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane2_r134 = 32'b100110_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane3_r134 = 32'b100110_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane4_r134 = 32'b100110_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane5_r134 = 32'b100110_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane6_r134 = 32'b100110_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane7_r134 = 32'b100110_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane8_r134 = 32'b100110_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane9_r134 = 32'b100110_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane10_r134 = 32'b100110_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane11_r134 = 32'b100110_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane12_r134 = 32'b100110_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane13_r134 = 32'b100110_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane14_r134 = 32'b100110_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane15_r134 = 32'b100110_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane16_r134 = 32'b100110_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane17_r134 = 32'b100110_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane18_r134 = 32'b100110_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane19_r134 = 32'b100110_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane20_r134 = 32'b100110_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane21_r134 = 32'b100110_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane22_r134 = 32'b100110_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane23_r134 = 32'b100110_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane24_r134 = 32'b100110_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane25_r134 = 32'b100110_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane26_r134 = 32'b100110_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane27_r134 = 32'b100110_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane28_r134 = 32'b100110_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane29_r134 = 32'b100110_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane30_r134 = 32'b100110_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.lane31_r134 = 32'b100110_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[38].pe.lane0_r135 = 32'b100110_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane1_r135 = 32'b100110_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane2_r135 = 32'b100110_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane3_r135 = 32'b100110_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane4_r135 = 32'b100110_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane5_r135 = 32'b100110_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane6_r135 = 32'b100110_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane7_r135 = 32'b100110_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane8_r135 = 32'b100110_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane9_r135 = 32'b100110_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane10_r135 = 32'b100110_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane11_r135 = 32'b100110_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane12_r135 = 32'b100110_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane13_r135 = 32'b100110_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane14_r135 = 32'b100110_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane15_r135 = 32'b100110_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane16_r135 = 32'b100110_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane17_r135 = 32'b100110_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane18_r135 = 32'b100110_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane19_r135 = 32'b100110_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane20_r135 = 32'b100110_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane21_r135 = 32'b100110_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane22_r135 = 32'b100110_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane23_r135 = 32'b100110_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane24_r135 = 32'b100110_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane25_r135 = 32'b100110_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane26_r135 = 32'b100110_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane27_r135 = 32'b100110_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane28_r135 = 32'b100110_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane29_r135 = 32'b100110_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane30_r135 = 32'b100110_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.lane31_r135 = 32'b100110_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[39].pe.lane0_r134 = 32'b100111_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane1_r134 = 32'b100111_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane2_r134 = 32'b100111_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane3_r134 = 32'b100111_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane4_r134 = 32'b100111_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane5_r134 = 32'b100111_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane6_r134 = 32'b100111_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane7_r134 = 32'b100111_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane8_r134 = 32'b100111_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane9_r134 = 32'b100111_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane10_r134 = 32'b100111_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane11_r134 = 32'b100111_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane12_r134 = 32'b100111_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane13_r134 = 32'b100111_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane14_r134 = 32'b100111_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane15_r134 = 32'b100111_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane16_r134 = 32'b100111_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane17_r134 = 32'b100111_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane18_r134 = 32'b100111_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane19_r134 = 32'b100111_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane20_r134 = 32'b100111_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane21_r134 = 32'b100111_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane22_r134 = 32'b100111_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane23_r134 = 32'b100111_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane24_r134 = 32'b100111_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane25_r134 = 32'b100111_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane26_r134 = 32'b100111_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane27_r134 = 32'b100111_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane28_r134 = 32'b100111_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane29_r134 = 32'b100111_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane30_r134 = 32'b100111_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.lane31_r134 = 32'b100111_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[39].pe.lane0_r135 = 32'b100111_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane1_r135 = 32'b100111_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane2_r135 = 32'b100111_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane3_r135 = 32'b100111_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane4_r135 = 32'b100111_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane5_r135 = 32'b100111_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane6_r135 = 32'b100111_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane7_r135 = 32'b100111_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane8_r135 = 32'b100111_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane9_r135 = 32'b100111_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane10_r135 = 32'b100111_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane11_r135 = 32'b100111_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane12_r135 = 32'b100111_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane13_r135 = 32'b100111_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane14_r135 = 32'b100111_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane15_r135 = 32'b100111_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane16_r135 = 32'b100111_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane17_r135 = 32'b100111_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane18_r135 = 32'b100111_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane19_r135 = 32'b100111_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane20_r135 = 32'b100111_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane21_r135 = 32'b100111_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane22_r135 = 32'b100111_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane23_r135 = 32'b100111_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane24_r135 = 32'b100111_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane25_r135 = 32'b100111_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane26_r135 = 32'b100111_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane27_r135 = 32'b100111_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane28_r135 = 32'b100111_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane29_r135 = 32'b100111_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane30_r135 = 32'b100111_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.lane31_r135 = 32'b100111_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[40].pe.lane0_r134 = 32'b101000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane1_r134 = 32'b101000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane2_r134 = 32'b101000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane3_r134 = 32'b101000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane4_r134 = 32'b101000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane5_r134 = 32'b101000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane6_r134 = 32'b101000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane7_r134 = 32'b101000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane8_r134 = 32'b101000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane9_r134 = 32'b101000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane10_r134 = 32'b101000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane11_r134 = 32'b101000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane12_r134 = 32'b101000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane13_r134 = 32'b101000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane14_r134 = 32'b101000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane15_r134 = 32'b101000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane16_r134 = 32'b101000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane17_r134 = 32'b101000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane18_r134 = 32'b101000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane19_r134 = 32'b101000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane20_r134 = 32'b101000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane21_r134 = 32'b101000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane22_r134 = 32'b101000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane23_r134 = 32'b101000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane24_r134 = 32'b101000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane25_r134 = 32'b101000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane26_r134 = 32'b101000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane27_r134 = 32'b101000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane28_r134 = 32'b101000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane29_r134 = 32'b101000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane30_r134 = 32'b101000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.lane31_r134 = 32'b101000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[40].pe.lane0_r135 = 32'b101000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane1_r135 = 32'b101000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane2_r135 = 32'b101000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane3_r135 = 32'b101000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane4_r135 = 32'b101000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane5_r135 = 32'b101000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane6_r135 = 32'b101000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane7_r135 = 32'b101000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane8_r135 = 32'b101000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane9_r135 = 32'b101000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane10_r135 = 32'b101000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane11_r135 = 32'b101000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane12_r135 = 32'b101000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane13_r135 = 32'b101000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane14_r135 = 32'b101000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane15_r135 = 32'b101000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane16_r135 = 32'b101000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane17_r135 = 32'b101000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane18_r135 = 32'b101000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane19_r135 = 32'b101000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane20_r135 = 32'b101000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane21_r135 = 32'b101000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane22_r135 = 32'b101000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane23_r135 = 32'b101000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane24_r135 = 32'b101000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane25_r135 = 32'b101000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane26_r135 = 32'b101000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane27_r135 = 32'b101000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane28_r135 = 32'b101000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane29_r135 = 32'b101000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane30_r135 = 32'b101000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.lane31_r135 = 32'b101000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[41].pe.lane0_r134 = 32'b101001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane1_r134 = 32'b101001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane2_r134 = 32'b101001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane3_r134 = 32'b101001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane4_r134 = 32'b101001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane5_r134 = 32'b101001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane6_r134 = 32'b101001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane7_r134 = 32'b101001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane8_r134 = 32'b101001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane9_r134 = 32'b101001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane10_r134 = 32'b101001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane11_r134 = 32'b101001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane12_r134 = 32'b101001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane13_r134 = 32'b101001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane14_r134 = 32'b101001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane15_r134 = 32'b101001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane16_r134 = 32'b101001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane17_r134 = 32'b101001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane18_r134 = 32'b101001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane19_r134 = 32'b101001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane20_r134 = 32'b101001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane21_r134 = 32'b101001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane22_r134 = 32'b101001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane23_r134 = 32'b101001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane24_r134 = 32'b101001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane25_r134 = 32'b101001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane26_r134 = 32'b101001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane27_r134 = 32'b101001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane28_r134 = 32'b101001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane29_r134 = 32'b101001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane30_r134 = 32'b101001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.lane31_r134 = 32'b101001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[41].pe.lane0_r135 = 32'b101001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane1_r135 = 32'b101001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane2_r135 = 32'b101001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane3_r135 = 32'b101001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane4_r135 = 32'b101001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane5_r135 = 32'b101001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane6_r135 = 32'b101001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane7_r135 = 32'b101001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane8_r135 = 32'b101001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane9_r135 = 32'b101001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane10_r135 = 32'b101001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane11_r135 = 32'b101001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane12_r135 = 32'b101001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane13_r135 = 32'b101001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane14_r135 = 32'b101001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane15_r135 = 32'b101001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane16_r135 = 32'b101001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane17_r135 = 32'b101001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane18_r135 = 32'b101001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane19_r135 = 32'b101001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane20_r135 = 32'b101001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane21_r135 = 32'b101001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane22_r135 = 32'b101001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane23_r135 = 32'b101001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane24_r135 = 32'b101001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane25_r135 = 32'b101001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane26_r135 = 32'b101001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane27_r135 = 32'b101001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane28_r135 = 32'b101001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane29_r135 = 32'b101001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane30_r135 = 32'b101001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.lane31_r135 = 32'b101001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[42].pe.lane0_r134 = 32'b101010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane1_r134 = 32'b101010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane2_r134 = 32'b101010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane3_r134 = 32'b101010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane4_r134 = 32'b101010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane5_r134 = 32'b101010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane6_r134 = 32'b101010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane7_r134 = 32'b101010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane8_r134 = 32'b101010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane9_r134 = 32'b101010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane10_r134 = 32'b101010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane11_r134 = 32'b101010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane12_r134 = 32'b101010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane13_r134 = 32'b101010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane14_r134 = 32'b101010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane15_r134 = 32'b101010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane16_r134 = 32'b101010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane17_r134 = 32'b101010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane18_r134 = 32'b101010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane19_r134 = 32'b101010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane20_r134 = 32'b101010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane21_r134 = 32'b101010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane22_r134 = 32'b101010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane23_r134 = 32'b101010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane24_r134 = 32'b101010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane25_r134 = 32'b101010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane26_r134 = 32'b101010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane27_r134 = 32'b101010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane28_r134 = 32'b101010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane29_r134 = 32'b101010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane30_r134 = 32'b101010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.lane31_r134 = 32'b101010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[42].pe.lane0_r135 = 32'b101010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane1_r135 = 32'b101010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane2_r135 = 32'b101010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane3_r135 = 32'b101010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane4_r135 = 32'b101010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane5_r135 = 32'b101010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane6_r135 = 32'b101010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane7_r135 = 32'b101010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane8_r135 = 32'b101010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane9_r135 = 32'b101010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane10_r135 = 32'b101010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane11_r135 = 32'b101010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane12_r135 = 32'b101010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane13_r135 = 32'b101010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane14_r135 = 32'b101010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane15_r135 = 32'b101010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane16_r135 = 32'b101010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane17_r135 = 32'b101010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane18_r135 = 32'b101010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane19_r135 = 32'b101010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane20_r135 = 32'b101010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane21_r135 = 32'b101010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane22_r135 = 32'b101010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane23_r135 = 32'b101010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane24_r135 = 32'b101010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane25_r135 = 32'b101010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane26_r135 = 32'b101010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane27_r135 = 32'b101010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane28_r135 = 32'b101010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane29_r135 = 32'b101010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane30_r135 = 32'b101010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.lane31_r135 = 32'b101010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[43].pe.lane0_r134 = 32'b101011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane1_r134 = 32'b101011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane2_r134 = 32'b101011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane3_r134 = 32'b101011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane4_r134 = 32'b101011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane5_r134 = 32'b101011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane6_r134 = 32'b101011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane7_r134 = 32'b101011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane8_r134 = 32'b101011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane9_r134 = 32'b101011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane10_r134 = 32'b101011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane11_r134 = 32'b101011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane12_r134 = 32'b101011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane13_r134 = 32'b101011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane14_r134 = 32'b101011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane15_r134 = 32'b101011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane16_r134 = 32'b101011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane17_r134 = 32'b101011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane18_r134 = 32'b101011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane19_r134 = 32'b101011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane20_r134 = 32'b101011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane21_r134 = 32'b101011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane22_r134 = 32'b101011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane23_r134 = 32'b101011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane24_r134 = 32'b101011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane25_r134 = 32'b101011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane26_r134 = 32'b101011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane27_r134 = 32'b101011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane28_r134 = 32'b101011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane29_r134 = 32'b101011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane30_r134 = 32'b101011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.lane31_r134 = 32'b101011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[43].pe.lane0_r135 = 32'b101011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane1_r135 = 32'b101011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane2_r135 = 32'b101011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane3_r135 = 32'b101011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane4_r135 = 32'b101011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane5_r135 = 32'b101011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane6_r135 = 32'b101011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane7_r135 = 32'b101011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane8_r135 = 32'b101011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane9_r135 = 32'b101011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane10_r135 = 32'b101011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane11_r135 = 32'b101011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane12_r135 = 32'b101011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane13_r135 = 32'b101011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane14_r135 = 32'b101011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane15_r135 = 32'b101011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane16_r135 = 32'b101011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane17_r135 = 32'b101011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane18_r135 = 32'b101011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane19_r135 = 32'b101011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane20_r135 = 32'b101011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane21_r135 = 32'b101011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane22_r135 = 32'b101011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane23_r135 = 32'b101011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane24_r135 = 32'b101011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane25_r135 = 32'b101011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane26_r135 = 32'b101011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane27_r135 = 32'b101011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane28_r135 = 32'b101011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane29_r135 = 32'b101011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane30_r135 = 32'b101011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.lane31_r135 = 32'b101011_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[44].pe.lane0_r134 = 32'b101100_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane1_r134 = 32'b101100_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane2_r134 = 32'b101100_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane3_r134 = 32'b101100_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane4_r134 = 32'b101100_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane5_r134 = 32'b101100_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane6_r134 = 32'b101100_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane7_r134 = 32'b101100_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane8_r134 = 32'b101100_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane9_r134 = 32'b101100_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane10_r134 = 32'b101100_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane11_r134 = 32'b101100_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane12_r134 = 32'b101100_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane13_r134 = 32'b101100_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane14_r134 = 32'b101100_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane15_r134 = 32'b101100_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane16_r134 = 32'b101100_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane17_r134 = 32'b101100_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane18_r134 = 32'b101100_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane19_r134 = 32'b101100_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane20_r134 = 32'b101100_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane21_r134 = 32'b101100_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane22_r134 = 32'b101100_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane23_r134 = 32'b101100_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane24_r134 = 32'b101100_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane25_r134 = 32'b101100_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane26_r134 = 32'b101100_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane27_r134 = 32'b101100_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane28_r134 = 32'b101100_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane29_r134 = 32'b101100_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane30_r134 = 32'b101100_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.lane31_r134 = 32'b101100_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[44].pe.lane0_r135 = 32'b101100_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane1_r135 = 32'b101100_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane2_r135 = 32'b101100_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane3_r135 = 32'b101100_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane4_r135 = 32'b101100_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane5_r135 = 32'b101100_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane6_r135 = 32'b101100_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane7_r135 = 32'b101100_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane8_r135 = 32'b101100_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane9_r135 = 32'b101100_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane10_r135 = 32'b101100_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane11_r135 = 32'b101100_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane12_r135 = 32'b101100_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane13_r135 = 32'b101100_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane14_r135 = 32'b101100_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane15_r135 = 32'b101100_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane16_r135 = 32'b101100_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane17_r135 = 32'b101100_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane18_r135 = 32'b101100_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane19_r135 = 32'b101100_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane20_r135 = 32'b101100_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane21_r135 = 32'b101100_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane22_r135 = 32'b101100_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane23_r135 = 32'b101100_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane24_r135 = 32'b101100_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane25_r135 = 32'b101100_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane26_r135 = 32'b101100_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane27_r135 = 32'b101100_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane28_r135 = 32'b101100_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane29_r135 = 32'b101100_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane30_r135 = 32'b101100_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.lane31_r135 = 32'b101100_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[45].pe.lane0_r134 = 32'b101101_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane1_r134 = 32'b101101_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane2_r134 = 32'b101101_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane3_r134 = 32'b101101_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane4_r134 = 32'b101101_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane5_r134 = 32'b101101_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane6_r134 = 32'b101101_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane7_r134 = 32'b101101_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane8_r134 = 32'b101101_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane9_r134 = 32'b101101_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane10_r134 = 32'b101101_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane11_r134 = 32'b101101_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane12_r134 = 32'b101101_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane13_r134 = 32'b101101_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane14_r134 = 32'b101101_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane15_r134 = 32'b101101_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane16_r134 = 32'b101101_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane17_r134 = 32'b101101_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane18_r134 = 32'b101101_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane19_r134 = 32'b101101_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane20_r134 = 32'b101101_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane21_r134 = 32'b101101_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane22_r134 = 32'b101101_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane23_r134 = 32'b101101_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane24_r134 = 32'b101101_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane25_r134 = 32'b101101_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane26_r134 = 32'b101101_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane27_r134 = 32'b101101_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane28_r134 = 32'b101101_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane29_r134 = 32'b101101_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane30_r134 = 32'b101101_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.lane31_r134 = 32'b101101_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[45].pe.lane0_r135 = 32'b101101_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane1_r135 = 32'b101101_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane2_r135 = 32'b101101_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane3_r135 = 32'b101101_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane4_r135 = 32'b101101_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane5_r135 = 32'b101101_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane6_r135 = 32'b101101_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane7_r135 = 32'b101101_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane8_r135 = 32'b101101_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane9_r135 = 32'b101101_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane10_r135 = 32'b101101_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane11_r135 = 32'b101101_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane12_r135 = 32'b101101_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane13_r135 = 32'b101101_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane14_r135 = 32'b101101_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane15_r135 = 32'b101101_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane16_r135 = 32'b101101_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane17_r135 = 32'b101101_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane18_r135 = 32'b101101_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane19_r135 = 32'b101101_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane20_r135 = 32'b101101_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane21_r135 = 32'b101101_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane22_r135 = 32'b101101_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane23_r135 = 32'b101101_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane24_r135 = 32'b101101_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane25_r135 = 32'b101101_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane26_r135 = 32'b101101_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane27_r135 = 32'b101101_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane28_r135 = 32'b101101_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane29_r135 = 32'b101101_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane30_r135 = 32'b101101_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.lane31_r135 = 32'b101101_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[46].pe.lane0_r134 = 32'b101110_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane1_r134 = 32'b101110_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane2_r134 = 32'b101110_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane3_r134 = 32'b101110_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane4_r134 = 32'b101110_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane5_r134 = 32'b101110_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane6_r134 = 32'b101110_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane7_r134 = 32'b101110_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane8_r134 = 32'b101110_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane9_r134 = 32'b101110_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane10_r134 = 32'b101110_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane11_r134 = 32'b101110_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane12_r134 = 32'b101110_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane13_r134 = 32'b101110_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane14_r134 = 32'b101110_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane15_r134 = 32'b101110_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane16_r134 = 32'b101110_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane17_r134 = 32'b101110_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane18_r134 = 32'b101110_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane19_r134 = 32'b101110_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane20_r134 = 32'b101110_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane21_r134 = 32'b101110_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane22_r134 = 32'b101110_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane23_r134 = 32'b101110_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane24_r134 = 32'b101110_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane25_r134 = 32'b101110_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane26_r134 = 32'b101110_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane27_r134 = 32'b101110_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane28_r134 = 32'b101110_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane29_r134 = 32'b101110_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane30_r134 = 32'b101110_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.lane31_r134 = 32'b101110_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[46].pe.lane0_r135 = 32'b101110_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane1_r135 = 32'b101110_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane2_r135 = 32'b101110_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane3_r135 = 32'b101110_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane4_r135 = 32'b101110_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane5_r135 = 32'b101110_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane6_r135 = 32'b101110_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane7_r135 = 32'b101110_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane8_r135 = 32'b101110_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane9_r135 = 32'b101110_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane10_r135 = 32'b101110_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane11_r135 = 32'b101110_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane12_r135 = 32'b101110_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane13_r135 = 32'b101110_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane14_r135 = 32'b101110_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane15_r135 = 32'b101110_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane16_r135 = 32'b101110_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane17_r135 = 32'b101110_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane18_r135 = 32'b101110_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane19_r135 = 32'b101110_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane20_r135 = 32'b101110_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane21_r135 = 32'b101110_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane22_r135 = 32'b101110_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane23_r135 = 32'b101110_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane24_r135 = 32'b101110_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane25_r135 = 32'b101110_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane26_r135 = 32'b101110_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane27_r135 = 32'b101110_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane28_r135 = 32'b101110_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane29_r135 = 32'b101110_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane30_r135 = 32'b101110_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.lane31_r135 = 32'b101110_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[47].pe.lane0_r134 = 32'b101111_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane1_r134 = 32'b101111_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane2_r134 = 32'b101111_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane3_r134 = 32'b101111_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane4_r134 = 32'b101111_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane5_r134 = 32'b101111_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane6_r134 = 32'b101111_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane7_r134 = 32'b101111_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane8_r134 = 32'b101111_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane9_r134 = 32'b101111_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane10_r134 = 32'b101111_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane11_r134 = 32'b101111_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane12_r134 = 32'b101111_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane13_r134 = 32'b101111_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane14_r134 = 32'b101111_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane15_r134 = 32'b101111_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane16_r134 = 32'b101111_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane17_r134 = 32'b101111_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane18_r134 = 32'b101111_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane19_r134 = 32'b101111_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane20_r134 = 32'b101111_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane21_r134 = 32'b101111_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane22_r134 = 32'b101111_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane23_r134 = 32'b101111_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane24_r134 = 32'b101111_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane25_r134 = 32'b101111_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane26_r134 = 32'b101111_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane27_r134 = 32'b101111_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane28_r134 = 32'b101111_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane29_r134 = 32'b101111_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane30_r134 = 32'b101111_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.lane31_r134 = 32'b101111_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[47].pe.lane0_r135 = 32'b101111_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane1_r135 = 32'b101111_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane2_r135 = 32'b101111_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane3_r135 = 32'b101111_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane4_r135 = 32'b101111_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane5_r135 = 32'b101111_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane6_r135 = 32'b101111_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane7_r135 = 32'b101111_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane8_r135 = 32'b101111_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane9_r135 = 32'b101111_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane10_r135 = 32'b101111_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane11_r135 = 32'b101111_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane12_r135 = 32'b101111_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane13_r135 = 32'b101111_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane14_r135 = 32'b101111_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane15_r135 = 32'b101111_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane16_r135 = 32'b101111_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane17_r135 = 32'b101111_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane18_r135 = 32'b101111_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane19_r135 = 32'b101111_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane20_r135 = 32'b101111_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane21_r135 = 32'b101111_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane22_r135 = 32'b101111_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane23_r135 = 32'b101111_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane24_r135 = 32'b101111_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane25_r135 = 32'b101111_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane26_r135 = 32'b101111_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane27_r135 = 32'b101111_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane28_r135 = 32'b101111_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane29_r135 = 32'b101111_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane30_r135 = 32'b101111_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.lane31_r135 = 32'b101111_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[48].pe.lane0_r134 = 32'b110000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane1_r134 = 32'b110000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane2_r134 = 32'b110000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane3_r134 = 32'b110000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane4_r134 = 32'b110000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane5_r134 = 32'b110000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane6_r134 = 32'b110000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane7_r134 = 32'b110000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane8_r134 = 32'b110000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane9_r134 = 32'b110000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane10_r134 = 32'b110000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane11_r134 = 32'b110000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane12_r134 = 32'b110000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane13_r134 = 32'b110000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane14_r134 = 32'b110000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane15_r134 = 32'b110000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane16_r134 = 32'b110000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane17_r134 = 32'b110000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane18_r134 = 32'b110000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane19_r134 = 32'b110000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane20_r134 = 32'b110000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane21_r134 = 32'b110000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane22_r134 = 32'b110000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane23_r134 = 32'b110000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane24_r134 = 32'b110000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane25_r134 = 32'b110000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane26_r134 = 32'b110000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane27_r134 = 32'b110000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane28_r134 = 32'b110000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane29_r134 = 32'b110000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane30_r134 = 32'b110000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.lane31_r134 = 32'b110000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[48].pe.lane0_r135 = 32'b110000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane1_r135 = 32'b110000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane2_r135 = 32'b110000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane3_r135 = 32'b110000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane4_r135 = 32'b110000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane5_r135 = 32'b110000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane6_r135 = 32'b110000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane7_r135 = 32'b110000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane8_r135 = 32'b110000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane9_r135 = 32'b110000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane10_r135 = 32'b110000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane11_r135 = 32'b110000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane12_r135 = 32'b110000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane13_r135 = 32'b110000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane14_r135 = 32'b110000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane15_r135 = 32'b110000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane16_r135 = 32'b110000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane17_r135 = 32'b110000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane18_r135 = 32'b110000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane19_r135 = 32'b110000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane20_r135 = 32'b110000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane21_r135 = 32'b110000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane22_r135 = 32'b110000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane23_r135 = 32'b110000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane24_r135 = 32'b110000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane25_r135 = 32'b110000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane26_r135 = 32'b110000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane27_r135 = 32'b110000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane28_r135 = 32'b110000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane29_r135 = 32'b110000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane30_r135 = 32'b110000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.lane31_r135 = 32'b110000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[49].pe.lane0_r134 = 32'b110001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane1_r134 = 32'b110001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane2_r134 = 32'b110001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane3_r134 = 32'b110001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane4_r134 = 32'b110001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane5_r134 = 32'b110001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane6_r134 = 32'b110001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane7_r134 = 32'b110001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane8_r134 = 32'b110001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane9_r134 = 32'b110001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane10_r134 = 32'b110001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane11_r134 = 32'b110001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane12_r134 = 32'b110001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane13_r134 = 32'b110001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane14_r134 = 32'b110001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane15_r134 = 32'b110001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane16_r134 = 32'b110001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane17_r134 = 32'b110001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane18_r134 = 32'b110001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane19_r134 = 32'b110001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane20_r134 = 32'b110001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane21_r134 = 32'b110001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane22_r134 = 32'b110001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane23_r134 = 32'b110001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane24_r134 = 32'b110001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane25_r134 = 32'b110001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane26_r134 = 32'b110001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane27_r134 = 32'b110001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane28_r134 = 32'b110001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane29_r134 = 32'b110001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane30_r134 = 32'b110001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.lane31_r134 = 32'b110001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[49].pe.lane0_r135 = 32'b110001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane1_r135 = 32'b110001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane2_r135 = 32'b110001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane3_r135 = 32'b110001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane4_r135 = 32'b110001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane5_r135 = 32'b110001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane6_r135 = 32'b110001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane7_r135 = 32'b110001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane8_r135 = 32'b110001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane9_r135 = 32'b110001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane10_r135 = 32'b110001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane11_r135 = 32'b110001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane12_r135 = 32'b110001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane13_r135 = 32'b110001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane14_r135 = 32'b110001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane15_r135 = 32'b110001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane16_r135 = 32'b110001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane17_r135 = 32'b110001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane18_r135 = 32'b110001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane19_r135 = 32'b110001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane20_r135 = 32'b110001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane21_r135 = 32'b110001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane22_r135 = 32'b110001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane23_r135 = 32'b110001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane24_r135 = 32'b110001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane25_r135 = 32'b110001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane26_r135 = 32'b110001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane27_r135 = 32'b110001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane28_r135 = 32'b110001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane29_r135 = 32'b110001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane30_r135 = 32'b110001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.lane31_r135 = 32'b110001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[50].pe.lane0_r134 = 32'b110010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane1_r134 = 32'b110010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane2_r134 = 32'b110010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane3_r134 = 32'b110010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane4_r134 = 32'b110010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane5_r134 = 32'b110010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane6_r134 = 32'b110010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane7_r134 = 32'b110010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane8_r134 = 32'b110010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane9_r134 = 32'b110010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane10_r134 = 32'b110010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane11_r134 = 32'b110010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane12_r134 = 32'b110010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane13_r134 = 32'b110010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane14_r134 = 32'b110010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane15_r134 = 32'b110010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane16_r134 = 32'b110010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane17_r134 = 32'b110010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane18_r134 = 32'b110010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane19_r134 = 32'b110010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane20_r134 = 32'b110010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane21_r134 = 32'b110010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane22_r134 = 32'b110010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane23_r134 = 32'b110010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane24_r134 = 32'b110010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane25_r134 = 32'b110010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane26_r134 = 32'b110010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane27_r134 = 32'b110010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane28_r134 = 32'b110010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane29_r134 = 32'b110010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane30_r134 = 32'b110010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.lane31_r134 = 32'b110010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[50].pe.lane0_r135 = 32'b110010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane1_r135 = 32'b110010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane2_r135 = 32'b110010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane3_r135 = 32'b110010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane4_r135 = 32'b110010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane5_r135 = 32'b110010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane6_r135 = 32'b110010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane7_r135 = 32'b110010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane8_r135 = 32'b110010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane9_r135 = 32'b110010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane10_r135 = 32'b110010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane11_r135 = 32'b110010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane12_r135 = 32'b110010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane13_r135 = 32'b110010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane14_r135 = 32'b110010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane15_r135 = 32'b110010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane16_r135 = 32'b110010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane17_r135 = 32'b110010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane18_r135 = 32'b110010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane19_r135 = 32'b110010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane20_r135 = 32'b110010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane21_r135 = 32'b110010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane22_r135 = 32'b110010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane23_r135 = 32'b110010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane24_r135 = 32'b110010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane25_r135 = 32'b110010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane26_r135 = 32'b110010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane27_r135 = 32'b110010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane28_r135 = 32'b110010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane29_r135 = 32'b110010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane30_r135 = 32'b110010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.lane31_r135 = 32'b110010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[51].pe.lane0_r134 = 32'b110011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane1_r134 = 32'b110011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane2_r134 = 32'b110011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane3_r134 = 32'b110011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane4_r134 = 32'b110011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane5_r134 = 32'b110011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane6_r134 = 32'b110011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane7_r134 = 32'b110011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane8_r134 = 32'b110011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane9_r134 = 32'b110011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane10_r134 = 32'b110011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane11_r134 = 32'b110011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane12_r134 = 32'b110011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane13_r134 = 32'b110011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane14_r134 = 32'b110011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane15_r134 = 32'b110011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane16_r134 = 32'b110011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane17_r134 = 32'b110011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane18_r134 = 32'b110011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane19_r134 = 32'b110011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane20_r134 = 32'b110011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane21_r134 = 32'b110011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane22_r134 = 32'b110011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane23_r134 = 32'b110011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane24_r134 = 32'b110011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane25_r134 = 32'b110011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane26_r134 = 32'b110011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane27_r134 = 32'b110011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane28_r134 = 32'b110011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane29_r134 = 32'b110011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane30_r134 = 32'b110011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.lane31_r134 = 32'b110011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[51].pe.lane0_r135 = 32'b110011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane1_r135 = 32'b110011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane2_r135 = 32'b110011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane3_r135 = 32'b110011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane4_r135 = 32'b110011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane5_r135 = 32'b110011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane6_r135 = 32'b110011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane7_r135 = 32'b110011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane8_r135 = 32'b110011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane9_r135 = 32'b110011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane10_r135 = 32'b110011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane11_r135 = 32'b110011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane12_r135 = 32'b110011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane13_r135 = 32'b110011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane14_r135 = 32'b110011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane15_r135 = 32'b110011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane16_r135 = 32'b110011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane17_r135 = 32'b110011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane18_r135 = 32'b110011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane19_r135 = 32'b110011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane20_r135 = 32'b110011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane21_r135 = 32'b110011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane22_r135 = 32'b110011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane23_r135 = 32'b110011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane24_r135 = 32'b110011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane25_r135 = 32'b110011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane26_r135 = 32'b110011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane27_r135 = 32'b110011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane28_r135 = 32'b110011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane29_r135 = 32'b110011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane30_r135 = 32'b110011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.lane31_r135 = 32'b110011_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[52].pe.lane0_r134 = 32'b110100_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane1_r134 = 32'b110100_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane2_r134 = 32'b110100_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane3_r134 = 32'b110100_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane4_r134 = 32'b110100_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane5_r134 = 32'b110100_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane6_r134 = 32'b110100_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane7_r134 = 32'b110100_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane8_r134 = 32'b110100_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane9_r134 = 32'b110100_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane10_r134 = 32'b110100_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane11_r134 = 32'b110100_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane12_r134 = 32'b110100_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane13_r134 = 32'b110100_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane14_r134 = 32'b110100_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane15_r134 = 32'b110100_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane16_r134 = 32'b110100_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane17_r134 = 32'b110100_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane18_r134 = 32'b110100_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane19_r134 = 32'b110100_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane20_r134 = 32'b110100_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane21_r134 = 32'b110100_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane22_r134 = 32'b110100_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane23_r134 = 32'b110100_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane24_r134 = 32'b110100_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane25_r134 = 32'b110100_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane26_r134 = 32'b110100_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane27_r134 = 32'b110100_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane28_r134 = 32'b110100_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane29_r134 = 32'b110100_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane30_r134 = 32'b110100_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.lane31_r134 = 32'b110100_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[52].pe.lane0_r135 = 32'b110100_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane1_r135 = 32'b110100_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane2_r135 = 32'b110100_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane3_r135 = 32'b110100_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane4_r135 = 32'b110100_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane5_r135 = 32'b110100_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane6_r135 = 32'b110100_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane7_r135 = 32'b110100_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane8_r135 = 32'b110100_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane9_r135 = 32'b110100_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane10_r135 = 32'b110100_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane11_r135 = 32'b110100_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane12_r135 = 32'b110100_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane13_r135 = 32'b110100_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane14_r135 = 32'b110100_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane15_r135 = 32'b110100_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane16_r135 = 32'b110100_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane17_r135 = 32'b110100_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane18_r135 = 32'b110100_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane19_r135 = 32'b110100_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane20_r135 = 32'b110100_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane21_r135 = 32'b110100_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane22_r135 = 32'b110100_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane23_r135 = 32'b110100_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane24_r135 = 32'b110100_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane25_r135 = 32'b110100_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane26_r135 = 32'b110100_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane27_r135 = 32'b110100_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane28_r135 = 32'b110100_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane29_r135 = 32'b110100_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane30_r135 = 32'b110100_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.lane31_r135 = 32'b110100_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[53].pe.lane0_r134 = 32'b110101_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane1_r134 = 32'b110101_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane2_r134 = 32'b110101_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane3_r134 = 32'b110101_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane4_r134 = 32'b110101_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane5_r134 = 32'b110101_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane6_r134 = 32'b110101_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane7_r134 = 32'b110101_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane8_r134 = 32'b110101_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane9_r134 = 32'b110101_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane10_r134 = 32'b110101_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane11_r134 = 32'b110101_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane12_r134 = 32'b110101_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane13_r134 = 32'b110101_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane14_r134 = 32'b110101_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane15_r134 = 32'b110101_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane16_r134 = 32'b110101_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane17_r134 = 32'b110101_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane18_r134 = 32'b110101_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane19_r134 = 32'b110101_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane20_r134 = 32'b110101_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane21_r134 = 32'b110101_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane22_r134 = 32'b110101_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane23_r134 = 32'b110101_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane24_r134 = 32'b110101_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane25_r134 = 32'b110101_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane26_r134 = 32'b110101_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane27_r134 = 32'b110101_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane28_r134 = 32'b110101_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane29_r134 = 32'b110101_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane30_r134 = 32'b110101_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.lane31_r134 = 32'b110101_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[53].pe.lane0_r135 = 32'b110101_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane1_r135 = 32'b110101_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane2_r135 = 32'b110101_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane3_r135 = 32'b110101_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane4_r135 = 32'b110101_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane5_r135 = 32'b110101_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane6_r135 = 32'b110101_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane7_r135 = 32'b110101_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane8_r135 = 32'b110101_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane9_r135 = 32'b110101_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane10_r135 = 32'b110101_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane11_r135 = 32'b110101_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane12_r135 = 32'b110101_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane13_r135 = 32'b110101_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane14_r135 = 32'b110101_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane15_r135 = 32'b110101_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane16_r135 = 32'b110101_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane17_r135 = 32'b110101_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane18_r135 = 32'b110101_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane19_r135 = 32'b110101_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane20_r135 = 32'b110101_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane21_r135 = 32'b110101_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane22_r135 = 32'b110101_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane23_r135 = 32'b110101_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane24_r135 = 32'b110101_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane25_r135 = 32'b110101_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane26_r135 = 32'b110101_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane27_r135 = 32'b110101_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane28_r135 = 32'b110101_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane29_r135 = 32'b110101_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane30_r135 = 32'b110101_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.lane31_r135 = 32'b110101_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[54].pe.lane0_r134 = 32'b110110_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane1_r134 = 32'b110110_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane2_r134 = 32'b110110_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane3_r134 = 32'b110110_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane4_r134 = 32'b110110_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane5_r134 = 32'b110110_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane6_r134 = 32'b110110_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane7_r134 = 32'b110110_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane8_r134 = 32'b110110_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane9_r134 = 32'b110110_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane10_r134 = 32'b110110_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane11_r134 = 32'b110110_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane12_r134 = 32'b110110_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane13_r134 = 32'b110110_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane14_r134 = 32'b110110_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane15_r134 = 32'b110110_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane16_r134 = 32'b110110_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane17_r134 = 32'b110110_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane18_r134 = 32'b110110_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane19_r134 = 32'b110110_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane20_r134 = 32'b110110_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane21_r134 = 32'b110110_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane22_r134 = 32'b110110_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane23_r134 = 32'b110110_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane24_r134 = 32'b110110_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane25_r134 = 32'b110110_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane26_r134 = 32'b110110_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane27_r134 = 32'b110110_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane28_r134 = 32'b110110_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane29_r134 = 32'b110110_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane30_r134 = 32'b110110_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.lane31_r134 = 32'b110110_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[54].pe.lane0_r135 = 32'b110110_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane1_r135 = 32'b110110_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane2_r135 = 32'b110110_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane3_r135 = 32'b110110_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane4_r135 = 32'b110110_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane5_r135 = 32'b110110_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane6_r135 = 32'b110110_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane7_r135 = 32'b110110_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane8_r135 = 32'b110110_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane9_r135 = 32'b110110_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane10_r135 = 32'b110110_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane11_r135 = 32'b110110_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane12_r135 = 32'b110110_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane13_r135 = 32'b110110_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane14_r135 = 32'b110110_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane15_r135 = 32'b110110_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane16_r135 = 32'b110110_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane17_r135 = 32'b110110_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane18_r135 = 32'b110110_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane19_r135 = 32'b110110_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane20_r135 = 32'b110110_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane21_r135 = 32'b110110_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane22_r135 = 32'b110110_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane23_r135 = 32'b110110_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane24_r135 = 32'b110110_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane25_r135 = 32'b110110_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane26_r135 = 32'b110110_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane27_r135 = 32'b110110_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane28_r135 = 32'b110110_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane29_r135 = 32'b110110_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane30_r135 = 32'b110110_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.lane31_r135 = 32'b110110_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[55].pe.lane0_r134 = 32'b110111_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane1_r134 = 32'b110111_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane2_r134 = 32'b110111_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane3_r134 = 32'b110111_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane4_r134 = 32'b110111_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane5_r134 = 32'b110111_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane6_r134 = 32'b110111_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane7_r134 = 32'b110111_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane8_r134 = 32'b110111_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane9_r134 = 32'b110111_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane10_r134 = 32'b110111_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane11_r134 = 32'b110111_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane12_r134 = 32'b110111_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane13_r134 = 32'b110111_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane14_r134 = 32'b110111_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane15_r134 = 32'b110111_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane16_r134 = 32'b110111_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane17_r134 = 32'b110111_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane18_r134 = 32'b110111_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane19_r134 = 32'b110111_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane20_r134 = 32'b110111_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane21_r134 = 32'b110111_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane22_r134 = 32'b110111_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane23_r134 = 32'b110111_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane24_r134 = 32'b110111_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane25_r134 = 32'b110111_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane26_r134 = 32'b110111_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane27_r134 = 32'b110111_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane28_r134 = 32'b110111_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane29_r134 = 32'b110111_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane30_r134 = 32'b110111_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.lane31_r134 = 32'b110111_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[55].pe.lane0_r135 = 32'b110111_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane1_r135 = 32'b110111_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane2_r135 = 32'b110111_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane3_r135 = 32'b110111_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane4_r135 = 32'b110111_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane5_r135 = 32'b110111_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane6_r135 = 32'b110111_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane7_r135 = 32'b110111_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane8_r135 = 32'b110111_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane9_r135 = 32'b110111_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane10_r135 = 32'b110111_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane11_r135 = 32'b110111_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane12_r135 = 32'b110111_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane13_r135 = 32'b110111_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane14_r135 = 32'b110111_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane15_r135 = 32'b110111_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane16_r135 = 32'b110111_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane17_r135 = 32'b110111_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane18_r135 = 32'b110111_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane19_r135 = 32'b110111_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane20_r135 = 32'b110111_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane21_r135 = 32'b110111_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane22_r135 = 32'b110111_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane23_r135 = 32'b110111_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane24_r135 = 32'b110111_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane25_r135 = 32'b110111_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane26_r135 = 32'b110111_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane27_r135 = 32'b110111_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane28_r135 = 32'b110111_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane29_r135 = 32'b110111_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane30_r135 = 32'b110111_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.lane31_r135 = 32'b110111_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[56].pe.lane0_r134 = 32'b111000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane1_r134 = 32'b111000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane2_r134 = 32'b111000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane3_r134 = 32'b111000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane4_r134 = 32'b111000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane5_r134 = 32'b111000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane6_r134 = 32'b111000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane7_r134 = 32'b111000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane8_r134 = 32'b111000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane9_r134 = 32'b111000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane10_r134 = 32'b111000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane11_r134 = 32'b111000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane12_r134 = 32'b111000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane13_r134 = 32'b111000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane14_r134 = 32'b111000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane15_r134 = 32'b111000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane16_r134 = 32'b111000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane17_r134 = 32'b111000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane18_r134 = 32'b111000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane19_r134 = 32'b111000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane20_r134 = 32'b111000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane21_r134 = 32'b111000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane22_r134 = 32'b111000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane23_r134 = 32'b111000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane24_r134 = 32'b111000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane25_r134 = 32'b111000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane26_r134 = 32'b111000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane27_r134 = 32'b111000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane28_r134 = 32'b111000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane29_r134 = 32'b111000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane30_r134 = 32'b111000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.lane31_r134 = 32'b111000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[56].pe.lane0_r135 = 32'b111000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane1_r135 = 32'b111000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane2_r135 = 32'b111000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane3_r135 = 32'b111000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane4_r135 = 32'b111000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane5_r135 = 32'b111000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane6_r135 = 32'b111000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane7_r135 = 32'b111000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane8_r135 = 32'b111000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane9_r135 = 32'b111000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane10_r135 = 32'b111000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane11_r135 = 32'b111000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane12_r135 = 32'b111000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane13_r135 = 32'b111000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane14_r135 = 32'b111000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane15_r135 = 32'b111000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane16_r135 = 32'b111000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane17_r135 = 32'b111000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane18_r135 = 32'b111000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane19_r135 = 32'b111000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane20_r135 = 32'b111000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane21_r135 = 32'b111000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane22_r135 = 32'b111000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane23_r135 = 32'b111000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane24_r135 = 32'b111000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane25_r135 = 32'b111000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane26_r135 = 32'b111000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane27_r135 = 32'b111000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane28_r135 = 32'b111000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane29_r135 = 32'b111000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane30_r135 = 32'b111000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.lane31_r135 = 32'b111000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[57].pe.lane0_r134 = 32'b111001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane1_r134 = 32'b111001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane2_r134 = 32'b111001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane3_r134 = 32'b111001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane4_r134 = 32'b111001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane5_r134 = 32'b111001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane6_r134 = 32'b111001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane7_r134 = 32'b111001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane8_r134 = 32'b111001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane9_r134 = 32'b111001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane10_r134 = 32'b111001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane11_r134 = 32'b111001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane12_r134 = 32'b111001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane13_r134 = 32'b111001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane14_r134 = 32'b111001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane15_r134 = 32'b111001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane16_r134 = 32'b111001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane17_r134 = 32'b111001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane18_r134 = 32'b111001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane19_r134 = 32'b111001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane20_r134 = 32'b111001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane21_r134 = 32'b111001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane22_r134 = 32'b111001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane23_r134 = 32'b111001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane24_r134 = 32'b111001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane25_r134 = 32'b111001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane26_r134 = 32'b111001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane27_r134 = 32'b111001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane28_r134 = 32'b111001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane29_r134 = 32'b111001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane30_r134 = 32'b111001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.lane31_r134 = 32'b111001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[57].pe.lane0_r135 = 32'b111001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane1_r135 = 32'b111001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane2_r135 = 32'b111001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane3_r135 = 32'b111001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane4_r135 = 32'b111001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane5_r135 = 32'b111001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane6_r135 = 32'b111001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane7_r135 = 32'b111001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane8_r135 = 32'b111001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane9_r135 = 32'b111001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane10_r135 = 32'b111001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane11_r135 = 32'b111001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane12_r135 = 32'b111001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane13_r135 = 32'b111001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane14_r135 = 32'b111001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane15_r135 = 32'b111001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane16_r135 = 32'b111001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane17_r135 = 32'b111001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane18_r135 = 32'b111001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane19_r135 = 32'b111001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane20_r135 = 32'b111001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane21_r135 = 32'b111001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane22_r135 = 32'b111001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane23_r135 = 32'b111001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane24_r135 = 32'b111001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane25_r135 = 32'b111001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane26_r135 = 32'b111001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane27_r135 = 32'b111001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane28_r135 = 32'b111001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane29_r135 = 32'b111001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane30_r135 = 32'b111001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.lane31_r135 = 32'b111001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[58].pe.lane0_r134 = 32'b111010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane1_r134 = 32'b111010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane2_r134 = 32'b111010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane3_r134 = 32'b111010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane4_r134 = 32'b111010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane5_r134 = 32'b111010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane6_r134 = 32'b111010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane7_r134 = 32'b111010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane8_r134 = 32'b111010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane9_r134 = 32'b111010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane10_r134 = 32'b111010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane11_r134 = 32'b111010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane12_r134 = 32'b111010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane13_r134 = 32'b111010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane14_r134 = 32'b111010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane15_r134 = 32'b111010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane16_r134 = 32'b111010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane17_r134 = 32'b111010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane18_r134 = 32'b111010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane19_r134 = 32'b111010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane20_r134 = 32'b111010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane21_r134 = 32'b111010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane22_r134 = 32'b111010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane23_r134 = 32'b111010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane24_r134 = 32'b111010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane25_r134 = 32'b111010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane26_r134 = 32'b111010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane27_r134 = 32'b111010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane28_r134 = 32'b111010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane29_r134 = 32'b111010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane30_r134 = 32'b111010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.lane31_r134 = 32'b111010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[58].pe.lane0_r135 = 32'b111010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane1_r135 = 32'b111010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane2_r135 = 32'b111010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane3_r135 = 32'b111010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane4_r135 = 32'b111010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane5_r135 = 32'b111010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane6_r135 = 32'b111010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane7_r135 = 32'b111010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane8_r135 = 32'b111010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane9_r135 = 32'b111010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane10_r135 = 32'b111010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane11_r135 = 32'b111010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane12_r135 = 32'b111010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane13_r135 = 32'b111010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane14_r135 = 32'b111010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane15_r135 = 32'b111010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane16_r135 = 32'b111010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane17_r135 = 32'b111010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane18_r135 = 32'b111010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane19_r135 = 32'b111010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane20_r135 = 32'b111010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane21_r135 = 32'b111010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane22_r135 = 32'b111010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane23_r135 = 32'b111010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane24_r135 = 32'b111010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane25_r135 = 32'b111010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane26_r135 = 32'b111010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane27_r135 = 32'b111010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane28_r135 = 32'b111010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane29_r135 = 32'b111010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane30_r135 = 32'b111010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.lane31_r135 = 32'b111010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[59].pe.lane0_r134 = 32'b111011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane1_r134 = 32'b111011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane2_r134 = 32'b111011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane3_r134 = 32'b111011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane4_r134 = 32'b111011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane5_r134 = 32'b111011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane6_r134 = 32'b111011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane7_r134 = 32'b111011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane8_r134 = 32'b111011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane9_r134 = 32'b111011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane10_r134 = 32'b111011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane11_r134 = 32'b111011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane12_r134 = 32'b111011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane13_r134 = 32'b111011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane14_r134 = 32'b111011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane15_r134 = 32'b111011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane16_r134 = 32'b111011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane17_r134 = 32'b111011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane18_r134 = 32'b111011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane19_r134 = 32'b111011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane20_r134 = 32'b111011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane21_r134 = 32'b111011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane22_r134 = 32'b111011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane23_r134 = 32'b111011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane24_r134 = 32'b111011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane25_r134 = 32'b111011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane26_r134 = 32'b111011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane27_r134 = 32'b111011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane28_r134 = 32'b111011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane29_r134 = 32'b111011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane30_r134 = 32'b111011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.lane31_r134 = 32'b111011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[59].pe.lane0_r135 = 32'b111011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane1_r135 = 32'b111011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane2_r135 = 32'b111011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane3_r135 = 32'b111011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane4_r135 = 32'b111011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane5_r135 = 32'b111011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane6_r135 = 32'b111011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane7_r135 = 32'b111011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane8_r135 = 32'b111011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane9_r135 = 32'b111011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane10_r135 = 32'b111011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane11_r135 = 32'b111011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane12_r135 = 32'b111011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane13_r135 = 32'b111011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane14_r135 = 32'b111011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane15_r135 = 32'b111011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane16_r135 = 32'b111011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane17_r135 = 32'b111011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane18_r135 = 32'b111011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane19_r135 = 32'b111011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane20_r135 = 32'b111011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane21_r135 = 32'b111011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane22_r135 = 32'b111011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane23_r135 = 32'b111011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane24_r135 = 32'b111011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane25_r135 = 32'b111011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane26_r135 = 32'b111011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane27_r135 = 32'b111011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane28_r135 = 32'b111011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane29_r135 = 32'b111011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane30_r135 = 32'b111011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.lane31_r135 = 32'b111011_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[60].pe.lane0_r134 = 32'b111100_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane1_r134 = 32'b111100_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane2_r134 = 32'b111100_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane3_r134 = 32'b111100_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane4_r134 = 32'b111100_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane5_r134 = 32'b111100_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane6_r134 = 32'b111100_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane7_r134 = 32'b111100_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane8_r134 = 32'b111100_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane9_r134 = 32'b111100_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane10_r134 = 32'b111100_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane11_r134 = 32'b111100_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane12_r134 = 32'b111100_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane13_r134 = 32'b111100_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane14_r134 = 32'b111100_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane15_r134 = 32'b111100_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane16_r134 = 32'b111100_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane17_r134 = 32'b111100_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane18_r134 = 32'b111100_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane19_r134 = 32'b111100_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane20_r134 = 32'b111100_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane21_r134 = 32'b111100_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane22_r134 = 32'b111100_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane23_r134 = 32'b111100_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane24_r134 = 32'b111100_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane25_r134 = 32'b111100_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane26_r134 = 32'b111100_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane27_r134 = 32'b111100_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane28_r134 = 32'b111100_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane29_r134 = 32'b111100_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane30_r134 = 32'b111100_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.lane31_r134 = 32'b111100_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[60].pe.lane0_r135 = 32'b111100_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane1_r135 = 32'b111100_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane2_r135 = 32'b111100_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane3_r135 = 32'b111100_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane4_r135 = 32'b111100_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane5_r135 = 32'b111100_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane6_r135 = 32'b111100_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane7_r135 = 32'b111100_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane8_r135 = 32'b111100_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane9_r135 = 32'b111100_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane10_r135 = 32'b111100_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane11_r135 = 32'b111100_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane12_r135 = 32'b111100_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane13_r135 = 32'b111100_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane14_r135 = 32'b111100_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane15_r135 = 32'b111100_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane16_r135 = 32'b111100_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane17_r135 = 32'b111100_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane18_r135 = 32'b111100_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane19_r135 = 32'b111100_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane20_r135 = 32'b111100_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane21_r135 = 32'b111100_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane22_r135 = 32'b111100_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane23_r135 = 32'b111100_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane24_r135 = 32'b111100_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane25_r135 = 32'b111100_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane26_r135 = 32'b111100_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane27_r135 = 32'b111100_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane28_r135 = 32'b111100_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane29_r135 = 32'b111100_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane30_r135 = 32'b111100_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.lane31_r135 = 32'b111100_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[61].pe.lane0_r134 = 32'b111101_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane1_r134 = 32'b111101_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane2_r134 = 32'b111101_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane3_r134 = 32'b111101_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane4_r134 = 32'b111101_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane5_r134 = 32'b111101_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane6_r134 = 32'b111101_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane7_r134 = 32'b111101_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane8_r134 = 32'b111101_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane9_r134 = 32'b111101_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane10_r134 = 32'b111101_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane11_r134 = 32'b111101_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane12_r134 = 32'b111101_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane13_r134 = 32'b111101_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane14_r134 = 32'b111101_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane15_r134 = 32'b111101_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane16_r134 = 32'b111101_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane17_r134 = 32'b111101_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane18_r134 = 32'b111101_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane19_r134 = 32'b111101_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane20_r134 = 32'b111101_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane21_r134 = 32'b111101_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane22_r134 = 32'b111101_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane23_r134 = 32'b111101_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane24_r134 = 32'b111101_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane25_r134 = 32'b111101_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane26_r134 = 32'b111101_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane27_r134 = 32'b111101_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane28_r134 = 32'b111101_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane29_r134 = 32'b111101_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane30_r134 = 32'b111101_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.lane31_r134 = 32'b111101_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[61].pe.lane0_r135 = 32'b111101_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane1_r135 = 32'b111101_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane2_r135 = 32'b111101_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane3_r135 = 32'b111101_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane4_r135 = 32'b111101_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane5_r135 = 32'b111101_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane6_r135 = 32'b111101_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane7_r135 = 32'b111101_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane8_r135 = 32'b111101_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane9_r135 = 32'b111101_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane10_r135 = 32'b111101_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane11_r135 = 32'b111101_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane12_r135 = 32'b111101_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane13_r135 = 32'b111101_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane14_r135 = 32'b111101_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane15_r135 = 32'b111101_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane16_r135 = 32'b111101_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane17_r135 = 32'b111101_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane18_r135 = 32'b111101_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane19_r135 = 32'b111101_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane20_r135 = 32'b111101_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane21_r135 = 32'b111101_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane22_r135 = 32'b111101_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane23_r135 = 32'b111101_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane24_r135 = 32'b111101_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane25_r135 = 32'b111101_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane26_r135 = 32'b111101_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane27_r135 = 32'b111101_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane28_r135 = 32'b111101_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane29_r135 = 32'b111101_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane30_r135 = 32'b111101_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.lane31_r135 = 32'b111101_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[62].pe.lane0_r134 = 32'b111110_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane1_r134 = 32'b111110_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane2_r134 = 32'b111110_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane3_r134 = 32'b111110_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane4_r134 = 32'b111110_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane5_r134 = 32'b111110_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane6_r134 = 32'b111110_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane7_r134 = 32'b111110_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane8_r134 = 32'b111110_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane9_r134 = 32'b111110_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane10_r134 = 32'b111110_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane11_r134 = 32'b111110_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane12_r134 = 32'b111110_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane13_r134 = 32'b111110_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane14_r134 = 32'b111110_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane15_r134 = 32'b111110_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane16_r134 = 32'b111110_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane17_r134 = 32'b111110_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane18_r134 = 32'b111110_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane19_r134 = 32'b111110_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane20_r134 = 32'b111110_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane21_r134 = 32'b111110_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane22_r134 = 32'b111110_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane23_r134 = 32'b111110_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane24_r134 = 32'b111110_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane25_r134 = 32'b111110_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane26_r134 = 32'b111110_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane27_r134 = 32'b111110_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane28_r134 = 32'b111110_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane29_r134 = 32'b111110_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane30_r134 = 32'b111110_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.lane31_r134 = 32'b111110_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[62].pe.lane0_r135 = 32'b111110_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane1_r135 = 32'b111110_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane2_r135 = 32'b111110_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane3_r135 = 32'b111110_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane4_r135 = 32'b111110_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane5_r135 = 32'b111110_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane6_r135 = 32'b111110_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane7_r135 = 32'b111110_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane8_r135 = 32'b111110_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane9_r135 = 32'b111110_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane10_r135 = 32'b111110_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane11_r135 = 32'b111110_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane12_r135 = 32'b111110_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane13_r135 = 32'b111110_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane14_r135 = 32'b111110_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane15_r135 = 32'b111110_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane16_r135 = 32'b111110_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane17_r135 = 32'b111110_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane18_r135 = 32'b111110_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane19_r135 = 32'b111110_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane20_r135 = 32'b111110_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane21_r135 = 32'b111110_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane22_r135 = 32'b111110_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane23_r135 = 32'b111110_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane24_r135 = 32'b111110_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane25_r135 = 32'b111110_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane26_r135 = 32'b111110_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane27_r135 = 32'b111110_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane28_r135 = 32'b111110_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane29_r135 = 32'b111110_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane30_r135 = 32'b111110_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.lane31_r135 = 32'b111110_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[63].pe.lane0_r134 = 32'b111111_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane1_r134 = 32'b111111_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane2_r134 = 32'b111111_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane3_r134 = 32'b111111_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane4_r134 = 32'b111111_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane5_r134 = 32'b111111_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane6_r134 = 32'b111111_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane7_r134 = 32'b111111_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane8_r134 = 32'b111111_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane9_r134 = 32'b111111_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane10_r134 = 32'b111111_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane11_r134 = 32'b111111_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane12_r134 = 32'b111111_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane13_r134 = 32'b111111_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane14_r134 = 32'b111111_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane15_r134 = 32'b111111_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane16_r134 = 32'b111111_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane17_r134 = 32'b111111_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane18_r134 = 32'b111111_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane19_r134 = 32'b111111_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane20_r134 = 32'b111111_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane21_r134 = 32'b111111_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane22_r134 = 32'b111111_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane23_r134 = 32'b111111_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane24_r134 = 32'b111111_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane25_r134 = 32'b111111_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane26_r134 = 32'b111111_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane27_r134 = 32'b111111_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane28_r134 = 32'b111111_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane29_r134 = 32'b111111_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane30_r134 = 32'b111111_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.lane31_r134 = 32'b111111_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[63].pe.lane0_r135 = 32'b111111_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane1_r135 = 32'b111111_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane2_r135 = 32'b111111_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane3_r135 = 32'b111111_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane4_r135 = 32'b111111_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane5_r135 = 32'b111111_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane6_r135 = 32'b111111_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane7_r135 = 32'b111111_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane8_r135 = 32'b111111_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane9_r135 = 32'b111111_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane10_r135 = 32'b111111_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane11_r135 = 32'b111111_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane12_r135 = 32'b111111_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane13_r135 = 32'b111111_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane14_r135 = 32'b111111_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane15_r135 = 32'b111111_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane16_r135 = 32'b111111_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane17_r135 = 32'b111111_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane18_r135 = 32'b111111_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane19_r135 = 32'b111111_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane20_r135 = 32'b111111_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane21_r135 = 32'b111111_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane22_r135 = 32'b111111_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane23_r135 = 32'b111111_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane24_r135 = 32'b111111_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane25_r135 = 32'b111111_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane26_r135 = 32'b111111_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane27_r135 = 32'b111111_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane28_r135 = 32'b111111_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane29_r135 = 32'b111111_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane30_r135 = 32'b111111_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.lane31_r135 = 32'b111111_11111__0_1000_0000_0000;

            // ##################################################
            // DMA Type and length of stream

            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[0].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[0].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[1].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[1].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[2].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[2].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[3].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[3].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[4].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[4].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[5].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[5].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[6].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[6].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[7].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[7].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[8].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[8].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[9].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[9].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[10].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[10].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[11].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[11].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[12].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[12].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[13].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[13].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[14].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[14].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[15].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[15].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[16].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[16].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[17].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[17].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[18].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[18].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[19].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[19].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[20].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[20].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[21].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[21].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[22].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[22].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[23].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[23].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[24].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[24].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[25].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[25].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[26].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[26].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[27].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[27].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[28].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[28].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[29].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[29].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[30].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[30].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[31].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[31].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[32].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[32].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[33].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[33].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[34].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[34].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[35].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[35].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[36].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[36].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[37].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[37].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[38].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[38].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[39].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[39].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[40].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[40].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[41].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[41].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[42].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[42].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[43].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[43].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[44].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[44].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[45].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[45].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[46].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[46].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[47].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[47].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[48].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[48].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[49].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[49].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[50].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[50].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[51].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[51].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[52].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[52].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[53].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[53].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[54].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[54].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[55].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[55].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[56].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[56].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[57].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[57].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[58].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[58].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[59].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[59].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[60].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[60].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[61].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[61].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[62].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[62].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[63].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[63].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane31_r133[15:0]  = numOfTypes;

            // ##################################################
            // Enable Stack bus streams

            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          
            enable_std_stream0 = 1 ;          
            enable_std_stream1 = 0 ;          

            // ##################################################
            // Enable and set transfer type

            repeat(10) @(negedge clk); 

            // Enable
            force pe_array_inst.pe_inst[0].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[1].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[2].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[3].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[4].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[5].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[6].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[7].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[8].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[9].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[10].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[11].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[12].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[13].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[14].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[15].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[16].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[17].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[18].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[19].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[20].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[21].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[22].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[23].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[24].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[25].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[26].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[27].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[28].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[29].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[30].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[31].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[32].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[33].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[34].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[35].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[36].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[37].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[38].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[39].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[40].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[41].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[42].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[43].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[44].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[45].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[46].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[47].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[48].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[49].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[50].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[51].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[52].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[53].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[54].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[55].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[56].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[57].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[58].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[59].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[60].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[61].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[62].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[63].pe.rs0[0]           = 1'b1;

            // Operation
            force pe_array_inst.pe_inst[0].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[1].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[2].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[3].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[4].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[5].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[6].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[7].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[8].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[9].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[10].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[11].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[12].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[13].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[14].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[15].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[16].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[17].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[18].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[19].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[20].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[21].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[22].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[23].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[24].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[25].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[26].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[27].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[28].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[29].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[30].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[31].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[32].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[33].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[34].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[35].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[36].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[37].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[38].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[39].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[40].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[41].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[42].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[43].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[44].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[45].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[46].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[47].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[48].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[49].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[50].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[51].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[52].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[53].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[54].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[55].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[56].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[57].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[58].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[59].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[60].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[61].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[62].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;
            force pe_array_inst.pe_inst[63].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM ;

            repeat(50) @(negedge clk);