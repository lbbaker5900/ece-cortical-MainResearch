
            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr0__std__oob_cntl                         ( mgr0__std__oob_cntl   ),
            .mgr0__std__oob_valid                        ( mgr0__std__oob_valid  ),
            .std__mgr0__oob_ready                        ( std__mgr0__oob_ready  ),
            .mgr0__std__oob_type                         ( mgr0__std__oob_type   ),
            .mgr0__std__oob_data                         ( mgr0__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr1__std__oob_cntl                         ( mgr1__std__oob_cntl   ),
            .mgr1__std__oob_valid                        ( mgr1__std__oob_valid  ),
            .std__mgr1__oob_ready                        ( std__mgr1__oob_ready  ),
            .mgr1__std__oob_type                         ( mgr1__std__oob_type   ),
            .mgr1__std__oob_data                         ( mgr1__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr2__std__oob_cntl                         ( mgr2__std__oob_cntl   ),
            .mgr2__std__oob_valid                        ( mgr2__std__oob_valid  ),
            .std__mgr2__oob_ready                        ( std__mgr2__oob_ready  ),
            .mgr2__std__oob_type                         ( mgr2__std__oob_type   ),
            .mgr2__std__oob_data                         ( mgr2__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr3__std__oob_cntl                         ( mgr3__std__oob_cntl   ),
            .mgr3__std__oob_valid                        ( mgr3__std__oob_valid  ),
            .std__mgr3__oob_ready                        ( std__mgr3__oob_ready  ),
            .mgr3__std__oob_type                         ( mgr3__std__oob_type   ),
            .mgr3__std__oob_data                         ( mgr3__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr4__std__oob_cntl                         ( mgr4__std__oob_cntl   ),
            .mgr4__std__oob_valid                        ( mgr4__std__oob_valid  ),
            .std__mgr4__oob_ready                        ( std__mgr4__oob_ready  ),
            .mgr4__std__oob_type                         ( mgr4__std__oob_type   ),
            .mgr4__std__oob_data                         ( mgr4__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr5__std__oob_cntl                         ( mgr5__std__oob_cntl   ),
            .mgr5__std__oob_valid                        ( mgr5__std__oob_valid  ),
            .std__mgr5__oob_ready                        ( std__mgr5__oob_ready  ),
            .mgr5__std__oob_type                         ( mgr5__std__oob_type   ),
            .mgr5__std__oob_data                         ( mgr5__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr6__std__oob_cntl                         ( mgr6__std__oob_cntl   ),
            .mgr6__std__oob_valid                        ( mgr6__std__oob_valid  ),
            .std__mgr6__oob_ready                        ( std__mgr6__oob_ready  ),
            .mgr6__std__oob_type                         ( mgr6__std__oob_type   ),
            .mgr6__std__oob_data                         ( mgr6__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr7__std__oob_cntl                         ( mgr7__std__oob_cntl   ),
            .mgr7__std__oob_valid                        ( mgr7__std__oob_valid  ),
            .std__mgr7__oob_ready                        ( std__mgr7__oob_ready  ),
            .mgr7__std__oob_type                         ( mgr7__std__oob_type   ),
            .mgr7__std__oob_data                         ( mgr7__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr8__std__oob_cntl                         ( mgr8__std__oob_cntl   ),
            .mgr8__std__oob_valid                        ( mgr8__std__oob_valid  ),
            .std__mgr8__oob_ready                        ( std__mgr8__oob_ready  ),
            .mgr8__std__oob_type                         ( mgr8__std__oob_type   ),
            .mgr8__std__oob_data                         ( mgr8__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr9__std__oob_cntl                         ( mgr9__std__oob_cntl   ),
            .mgr9__std__oob_valid                        ( mgr9__std__oob_valid  ),
            .std__mgr9__oob_ready                        ( std__mgr9__oob_ready  ),
            .mgr9__std__oob_type                         ( mgr9__std__oob_type   ),
            .mgr9__std__oob_data                         ( mgr9__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr10__std__oob_cntl                         ( mgr10__std__oob_cntl   ),
            .mgr10__std__oob_valid                        ( mgr10__std__oob_valid  ),
            .std__mgr10__oob_ready                        ( std__mgr10__oob_ready  ),
            .mgr10__std__oob_type                         ( mgr10__std__oob_type   ),
            .mgr10__std__oob_data                         ( mgr10__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr11__std__oob_cntl                         ( mgr11__std__oob_cntl   ),
            .mgr11__std__oob_valid                        ( mgr11__std__oob_valid  ),
            .std__mgr11__oob_ready                        ( std__mgr11__oob_ready  ),
            .mgr11__std__oob_type                         ( mgr11__std__oob_type   ),
            .mgr11__std__oob_data                         ( mgr11__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr12__std__oob_cntl                         ( mgr12__std__oob_cntl   ),
            .mgr12__std__oob_valid                        ( mgr12__std__oob_valid  ),
            .std__mgr12__oob_ready                        ( std__mgr12__oob_ready  ),
            .mgr12__std__oob_type                         ( mgr12__std__oob_type   ),
            .mgr12__std__oob_data                         ( mgr12__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr13__std__oob_cntl                         ( mgr13__std__oob_cntl   ),
            .mgr13__std__oob_valid                        ( mgr13__std__oob_valid  ),
            .std__mgr13__oob_ready                        ( std__mgr13__oob_ready  ),
            .mgr13__std__oob_type                         ( mgr13__std__oob_type   ),
            .mgr13__std__oob_data                         ( mgr13__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr14__std__oob_cntl                         ( mgr14__std__oob_cntl   ),
            .mgr14__std__oob_valid                        ( mgr14__std__oob_valid  ),
            .std__mgr14__oob_ready                        ( std__mgr14__oob_ready  ),
            .mgr14__std__oob_type                         ( mgr14__std__oob_type   ),
            .mgr14__std__oob_data                         ( mgr14__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr15__std__oob_cntl                         ( mgr15__std__oob_cntl   ),
            .mgr15__std__oob_valid                        ( mgr15__std__oob_valid  ),
            .std__mgr15__oob_ready                        ( std__mgr15__oob_ready  ),
            .mgr15__std__oob_type                         ( mgr15__std__oob_type   ),
            .mgr15__std__oob_data                         ( mgr15__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr16__std__oob_cntl                         ( mgr16__std__oob_cntl   ),
            .mgr16__std__oob_valid                        ( mgr16__std__oob_valid  ),
            .std__mgr16__oob_ready                        ( std__mgr16__oob_ready  ),
            .mgr16__std__oob_type                         ( mgr16__std__oob_type   ),
            .mgr16__std__oob_data                         ( mgr16__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr17__std__oob_cntl                         ( mgr17__std__oob_cntl   ),
            .mgr17__std__oob_valid                        ( mgr17__std__oob_valid  ),
            .std__mgr17__oob_ready                        ( std__mgr17__oob_ready  ),
            .mgr17__std__oob_type                         ( mgr17__std__oob_type   ),
            .mgr17__std__oob_data                         ( mgr17__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr18__std__oob_cntl                         ( mgr18__std__oob_cntl   ),
            .mgr18__std__oob_valid                        ( mgr18__std__oob_valid  ),
            .std__mgr18__oob_ready                        ( std__mgr18__oob_ready  ),
            .mgr18__std__oob_type                         ( mgr18__std__oob_type   ),
            .mgr18__std__oob_data                         ( mgr18__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr19__std__oob_cntl                         ( mgr19__std__oob_cntl   ),
            .mgr19__std__oob_valid                        ( mgr19__std__oob_valid  ),
            .std__mgr19__oob_ready                        ( std__mgr19__oob_ready  ),
            .mgr19__std__oob_type                         ( mgr19__std__oob_type   ),
            .mgr19__std__oob_data                         ( mgr19__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr20__std__oob_cntl                         ( mgr20__std__oob_cntl   ),
            .mgr20__std__oob_valid                        ( mgr20__std__oob_valid  ),
            .std__mgr20__oob_ready                        ( std__mgr20__oob_ready  ),
            .mgr20__std__oob_type                         ( mgr20__std__oob_type   ),
            .mgr20__std__oob_data                         ( mgr20__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr21__std__oob_cntl                         ( mgr21__std__oob_cntl   ),
            .mgr21__std__oob_valid                        ( mgr21__std__oob_valid  ),
            .std__mgr21__oob_ready                        ( std__mgr21__oob_ready  ),
            .mgr21__std__oob_type                         ( mgr21__std__oob_type   ),
            .mgr21__std__oob_data                         ( mgr21__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr22__std__oob_cntl                         ( mgr22__std__oob_cntl   ),
            .mgr22__std__oob_valid                        ( mgr22__std__oob_valid  ),
            .std__mgr22__oob_ready                        ( std__mgr22__oob_ready  ),
            .mgr22__std__oob_type                         ( mgr22__std__oob_type   ),
            .mgr22__std__oob_data                         ( mgr22__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr23__std__oob_cntl                         ( mgr23__std__oob_cntl   ),
            .mgr23__std__oob_valid                        ( mgr23__std__oob_valid  ),
            .std__mgr23__oob_ready                        ( std__mgr23__oob_ready  ),
            .mgr23__std__oob_type                         ( mgr23__std__oob_type   ),
            .mgr23__std__oob_data                         ( mgr23__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr24__std__oob_cntl                         ( mgr24__std__oob_cntl   ),
            .mgr24__std__oob_valid                        ( mgr24__std__oob_valid  ),
            .std__mgr24__oob_ready                        ( std__mgr24__oob_ready  ),
            .mgr24__std__oob_type                         ( mgr24__std__oob_type   ),
            .mgr24__std__oob_data                         ( mgr24__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr25__std__oob_cntl                         ( mgr25__std__oob_cntl   ),
            .mgr25__std__oob_valid                        ( mgr25__std__oob_valid  ),
            .std__mgr25__oob_ready                        ( std__mgr25__oob_ready  ),
            .mgr25__std__oob_type                         ( mgr25__std__oob_type   ),
            .mgr25__std__oob_data                         ( mgr25__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr26__std__oob_cntl                         ( mgr26__std__oob_cntl   ),
            .mgr26__std__oob_valid                        ( mgr26__std__oob_valid  ),
            .std__mgr26__oob_ready                        ( std__mgr26__oob_ready  ),
            .mgr26__std__oob_type                         ( mgr26__std__oob_type   ),
            .mgr26__std__oob_data                         ( mgr26__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr27__std__oob_cntl                         ( mgr27__std__oob_cntl   ),
            .mgr27__std__oob_valid                        ( mgr27__std__oob_valid  ),
            .std__mgr27__oob_ready                        ( std__mgr27__oob_ready  ),
            .mgr27__std__oob_type                         ( mgr27__std__oob_type   ),
            .mgr27__std__oob_data                         ( mgr27__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr28__std__oob_cntl                         ( mgr28__std__oob_cntl   ),
            .mgr28__std__oob_valid                        ( mgr28__std__oob_valid  ),
            .std__mgr28__oob_ready                        ( std__mgr28__oob_ready  ),
            .mgr28__std__oob_type                         ( mgr28__std__oob_type   ),
            .mgr28__std__oob_data                         ( mgr28__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr29__std__oob_cntl                         ( mgr29__std__oob_cntl   ),
            .mgr29__std__oob_valid                        ( mgr29__std__oob_valid  ),
            .std__mgr29__oob_ready                        ( std__mgr29__oob_ready  ),
            .mgr29__std__oob_type                         ( mgr29__std__oob_type   ),
            .mgr29__std__oob_data                         ( mgr29__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr30__std__oob_cntl                         ( mgr30__std__oob_cntl   ),
            .mgr30__std__oob_valid                        ( mgr30__std__oob_valid  ),
            .std__mgr30__oob_ready                        ( std__mgr30__oob_ready  ),
            .mgr30__std__oob_type                         ( mgr30__std__oob_type   ),
            .mgr30__std__oob_data                         ( mgr30__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr31__std__oob_cntl                         ( mgr31__std__oob_cntl   ),
            .mgr31__std__oob_valid                        ( mgr31__std__oob_valid  ),
            .std__mgr31__oob_ready                        ( std__mgr31__oob_ready  ),
            .mgr31__std__oob_type                         ( mgr31__std__oob_type   ),
            .mgr31__std__oob_data                         ( mgr31__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr32__std__oob_cntl                         ( mgr32__std__oob_cntl   ),
            .mgr32__std__oob_valid                        ( mgr32__std__oob_valid  ),
            .std__mgr32__oob_ready                        ( std__mgr32__oob_ready  ),
            .mgr32__std__oob_type                         ( mgr32__std__oob_type   ),
            .mgr32__std__oob_data                         ( mgr32__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr33__std__oob_cntl                         ( mgr33__std__oob_cntl   ),
            .mgr33__std__oob_valid                        ( mgr33__std__oob_valid  ),
            .std__mgr33__oob_ready                        ( std__mgr33__oob_ready  ),
            .mgr33__std__oob_type                         ( mgr33__std__oob_type   ),
            .mgr33__std__oob_data                         ( mgr33__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr34__std__oob_cntl                         ( mgr34__std__oob_cntl   ),
            .mgr34__std__oob_valid                        ( mgr34__std__oob_valid  ),
            .std__mgr34__oob_ready                        ( std__mgr34__oob_ready  ),
            .mgr34__std__oob_type                         ( mgr34__std__oob_type   ),
            .mgr34__std__oob_data                         ( mgr34__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr35__std__oob_cntl                         ( mgr35__std__oob_cntl   ),
            .mgr35__std__oob_valid                        ( mgr35__std__oob_valid  ),
            .std__mgr35__oob_ready                        ( std__mgr35__oob_ready  ),
            .mgr35__std__oob_type                         ( mgr35__std__oob_type   ),
            .mgr35__std__oob_data                         ( mgr35__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr36__std__oob_cntl                         ( mgr36__std__oob_cntl   ),
            .mgr36__std__oob_valid                        ( mgr36__std__oob_valid  ),
            .std__mgr36__oob_ready                        ( std__mgr36__oob_ready  ),
            .mgr36__std__oob_type                         ( mgr36__std__oob_type   ),
            .mgr36__std__oob_data                         ( mgr36__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr37__std__oob_cntl                         ( mgr37__std__oob_cntl   ),
            .mgr37__std__oob_valid                        ( mgr37__std__oob_valid  ),
            .std__mgr37__oob_ready                        ( std__mgr37__oob_ready  ),
            .mgr37__std__oob_type                         ( mgr37__std__oob_type   ),
            .mgr37__std__oob_data                         ( mgr37__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr38__std__oob_cntl                         ( mgr38__std__oob_cntl   ),
            .mgr38__std__oob_valid                        ( mgr38__std__oob_valid  ),
            .std__mgr38__oob_ready                        ( std__mgr38__oob_ready  ),
            .mgr38__std__oob_type                         ( mgr38__std__oob_type   ),
            .mgr38__std__oob_data                         ( mgr38__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr39__std__oob_cntl                         ( mgr39__std__oob_cntl   ),
            .mgr39__std__oob_valid                        ( mgr39__std__oob_valid  ),
            .std__mgr39__oob_ready                        ( std__mgr39__oob_ready  ),
            .mgr39__std__oob_type                         ( mgr39__std__oob_type   ),
            .mgr39__std__oob_data                         ( mgr39__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr40__std__oob_cntl                         ( mgr40__std__oob_cntl   ),
            .mgr40__std__oob_valid                        ( mgr40__std__oob_valid  ),
            .std__mgr40__oob_ready                        ( std__mgr40__oob_ready  ),
            .mgr40__std__oob_type                         ( mgr40__std__oob_type   ),
            .mgr40__std__oob_data                         ( mgr40__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr41__std__oob_cntl                         ( mgr41__std__oob_cntl   ),
            .mgr41__std__oob_valid                        ( mgr41__std__oob_valid  ),
            .std__mgr41__oob_ready                        ( std__mgr41__oob_ready  ),
            .mgr41__std__oob_type                         ( mgr41__std__oob_type   ),
            .mgr41__std__oob_data                         ( mgr41__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr42__std__oob_cntl                         ( mgr42__std__oob_cntl   ),
            .mgr42__std__oob_valid                        ( mgr42__std__oob_valid  ),
            .std__mgr42__oob_ready                        ( std__mgr42__oob_ready  ),
            .mgr42__std__oob_type                         ( mgr42__std__oob_type   ),
            .mgr42__std__oob_data                         ( mgr42__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr43__std__oob_cntl                         ( mgr43__std__oob_cntl   ),
            .mgr43__std__oob_valid                        ( mgr43__std__oob_valid  ),
            .std__mgr43__oob_ready                        ( std__mgr43__oob_ready  ),
            .mgr43__std__oob_type                         ( mgr43__std__oob_type   ),
            .mgr43__std__oob_data                         ( mgr43__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr44__std__oob_cntl                         ( mgr44__std__oob_cntl   ),
            .mgr44__std__oob_valid                        ( mgr44__std__oob_valid  ),
            .std__mgr44__oob_ready                        ( std__mgr44__oob_ready  ),
            .mgr44__std__oob_type                         ( mgr44__std__oob_type   ),
            .mgr44__std__oob_data                         ( mgr44__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr45__std__oob_cntl                         ( mgr45__std__oob_cntl   ),
            .mgr45__std__oob_valid                        ( mgr45__std__oob_valid  ),
            .std__mgr45__oob_ready                        ( std__mgr45__oob_ready  ),
            .mgr45__std__oob_type                         ( mgr45__std__oob_type   ),
            .mgr45__std__oob_data                         ( mgr45__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr46__std__oob_cntl                         ( mgr46__std__oob_cntl   ),
            .mgr46__std__oob_valid                        ( mgr46__std__oob_valid  ),
            .std__mgr46__oob_ready                        ( std__mgr46__oob_ready  ),
            .mgr46__std__oob_type                         ( mgr46__std__oob_type   ),
            .mgr46__std__oob_data                         ( mgr46__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr47__std__oob_cntl                         ( mgr47__std__oob_cntl   ),
            .mgr47__std__oob_valid                        ( mgr47__std__oob_valid  ),
            .std__mgr47__oob_ready                        ( std__mgr47__oob_ready  ),
            .mgr47__std__oob_type                         ( mgr47__std__oob_type   ),
            .mgr47__std__oob_data                         ( mgr47__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr48__std__oob_cntl                         ( mgr48__std__oob_cntl   ),
            .mgr48__std__oob_valid                        ( mgr48__std__oob_valid  ),
            .std__mgr48__oob_ready                        ( std__mgr48__oob_ready  ),
            .mgr48__std__oob_type                         ( mgr48__std__oob_type   ),
            .mgr48__std__oob_data                         ( mgr48__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr49__std__oob_cntl                         ( mgr49__std__oob_cntl   ),
            .mgr49__std__oob_valid                        ( mgr49__std__oob_valid  ),
            .std__mgr49__oob_ready                        ( std__mgr49__oob_ready  ),
            .mgr49__std__oob_type                         ( mgr49__std__oob_type   ),
            .mgr49__std__oob_data                         ( mgr49__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr50__std__oob_cntl                         ( mgr50__std__oob_cntl   ),
            .mgr50__std__oob_valid                        ( mgr50__std__oob_valid  ),
            .std__mgr50__oob_ready                        ( std__mgr50__oob_ready  ),
            .mgr50__std__oob_type                         ( mgr50__std__oob_type   ),
            .mgr50__std__oob_data                         ( mgr50__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr51__std__oob_cntl                         ( mgr51__std__oob_cntl   ),
            .mgr51__std__oob_valid                        ( mgr51__std__oob_valid  ),
            .std__mgr51__oob_ready                        ( std__mgr51__oob_ready  ),
            .mgr51__std__oob_type                         ( mgr51__std__oob_type   ),
            .mgr51__std__oob_data                         ( mgr51__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr52__std__oob_cntl                         ( mgr52__std__oob_cntl   ),
            .mgr52__std__oob_valid                        ( mgr52__std__oob_valid  ),
            .std__mgr52__oob_ready                        ( std__mgr52__oob_ready  ),
            .mgr52__std__oob_type                         ( mgr52__std__oob_type   ),
            .mgr52__std__oob_data                         ( mgr52__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr53__std__oob_cntl                         ( mgr53__std__oob_cntl   ),
            .mgr53__std__oob_valid                        ( mgr53__std__oob_valid  ),
            .std__mgr53__oob_ready                        ( std__mgr53__oob_ready  ),
            .mgr53__std__oob_type                         ( mgr53__std__oob_type   ),
            .mgr53__std__oob_data                         ( mgr53__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr54__std__oob_cntl                         ( mgr54__std__oob_cntl   ),
            .mgr54__std__oob_valid                        ( mgr54__std__oob_valid  ),
            .std__mgr54__oob_ready                        ( std__mgr54__oob_ready  ),
            .mgr54__std__oob_type                         ( mgr54__std__oob_type   ),
            .mgr54__std__oob_data                         ( mgr54__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr55__std__oob_cntl                         ( mgr55__std__oob_cntl   ),
            .mgr55__std__oob_valid                        ( mgr55__std__oob_valid  ),
            .std__mgr55__oob_ready                        ( std__mgr55__oob_ready  ),
            .mgr55__std__oob_type                         ( mgr55__std__oob_type   ),
            .mgr55__std__oob_data                         ( mgr55__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr56__std__oob_cntl                         ( mgr56__std__oob_cntl   ),
            .mgr56__std__oob_valid                        ( mgr56__std__oob_valid  ),
            .std__mgr56__oob_ready                        ( std__mgr56__oob_ready  ),
            .mgr56__std__oob_type                         ( mgr56__std__oob_type   ),
            .mgr56__std__oob_data                         ( mgr56__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr57__std__oob_cntl                         ( mgr57__std__oob_cntl   ),
            .mgr57__std__oob_valid                        ( mgr57__std__oob_valid  ),
            .std__mgr57__oob_ready                        ( std__mgr57__oob_ready  ),
            .mgr57__std__oob_type                         ( mgr57__std__oob_type   ),
            .mgr57__std__oob_data                         ( mgr57__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr58__std__oob_cntl                         ( mgr58__std__oob_cntl   ),
            .mgr58__std__oob_valid                        ( mgr58__std__oob_valid  ),
            .std__mgr58__oob_ready                        ( std__mgr58__oob_ready  ),
            .mgr58__std__oob_type                         ( mgr58__std__oob_type   ),
            .mgr58__std__oob_data                         ( mgr58__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr59__std__oob_cntl                         ( mgr59__std__oob_cntl   ),
            .mgr59__std__oob_valid                        ( mgr59__std__oob_valid  ),
            .std__mgr59__oob_ready                        ( std__mgr59__oob_ready  ),
            .mgr59__std__oob_type                         ( mgr59__std__oob_type   ),
            .mgr59__std__oob_data                         ( mgr59__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr60__std__oob_cntl                         ( mgr60__std__oob_cntl   ),
            .mgr60__std__oob_valid                        ( mgr60__std__oob_valid  ),
            .std__mgr60__oob_ready                        ( std__mgr60__oob_ready  ),
            .mgr60__std__oob_type                         ( mgr60__std__oob_type   ),
            .mgr60__std__oob_data                         ( mgr60__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr61__std__oob_cntl                         ( mgr61__std__oob_cntl   ),
            .mgr61__std__oob_valid                        ( mgr61__std__oob_valid  ),
            .std__mgr61__oob_ready                        ( std__mgr61__oob_ready  ),
            .mgr61__std__oob_type                         ( mgr61__std__oob_type   ),
            .mgr61__std__oob_data                         ( mgr61__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr62__std__oob_cntl                         ( mgr62__std__oob_cntl   ),
            .mgr62__std__oob_valid                        ( mgr62__std__oob_valid  ),
            .std__mgr62__oob_ready                        ( std__mgr62__oob_ready  ),
            .mgr62__std__oob_type                         ( mgr62__std__oob_type   ),
            .mgr62__std__oob_data                         ( mgr62__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr63__std__oob_cntl                         ( mgr63__std__oob_cntl   ),
            .mgr63__std__oob_valid                        ( mgr63__std__oob_valid  ),
            .std__mgr63__oob_ready                        ( std__mgr63__oob_ready  ),
            .mgr63__std__oob_type                         ( mgr63__std__oob_type   ),
            .mgr63__std__oob_data                         ( mgr63__std__oob_data   ),
