
  assign   rs0  = simd__scntl__rs0 ;
  assign   rs1  = simd__scntl__rs1 ;

// Lane 0                 
  assign   lane0_r128  =  simd__scntl__lane_r128 [0] ;
  assign   lane0_r129  =  simd__scntl__lane_r129 [0] ;
  assign   lane0_r130  =  simd__scntl__lane_r130 [0] ;
  assign   lane0_r131  =  simd__scntl__lane_r131 [0] ;
  assign   lane0_r132  =  simd__scntl__lane_r132 [0] ;
  assign   lane0_r133  =  simd__scntl__lane_r133 [0] ;
  assign   lane0_r134  =  simd__scntl__lane_r134 [0] ;
  assign   lane0_r135  =  simd__scntl__lane_r135 [0] ;

// Lane 1                 
  assign   lane1_r128  =  simd__scntl__lane_r128 [1] ;
  assign   lane1_r129  =  simd__scntl__lane_r129 [1] ;
  assign   lane1_r130  =  simd__scntl__lane_r130 [1] ;
  assign   lane1_r131  =  simd__scntl__lane_r131 [1] ;
  assign   lane1_r132  =  simd__scntl__lane_r132 [1] ;
  assign   lane1_r133  =  simd__scntl__lane_r133 [1] ;
  assign   lane1_r134  =  simd__scntl__lane_r134 [1] ;
  assign   lane1_r135  =  simd__scntl__lane_r135 [1] ;

// Lane 2                 
  assign   lane2_r128  =  simd__scntl__lane_r128 [2] ;
  assign   lane2_r129  =  simd__scntl__lane_r129 [2] ;
  assign   lane2_r130  =  simd__scntl__lane_r130 [2] ;
  assign   lane2_r131  =  simd__scntl__lane_r131 [2] ;
  assign   lane2_r132  =  simd__scntl__lane_r132 [2] ;
  assign   lane2_r133  =  simd__scntl__lane_r133 [2] ;
  assign   lane2_r134  =  simd__scntl__lane_r134 [2] ;
  assign   lane2_r135  =  simd__scntl__lane_r135 [2] ;

// Lane 3                 
  assign   lane3_r128  =  simd__scntl__lane_r128 [3] ;
  assign   lane3_r129  =  simd__scntl__lane_r129 [3] ;
  assign   lane3_r130  =  simd__scntl__lane_r130 [3] ;
  assign   lane3_r131  =  simd__scntl__lane_r131 [3] ;
  assign   lane3_r132  =  simd__scntl__lane_r132 [3] ;
  assign   lane3_r133  =  simd__scntl__lane_r133 [3] ;
  assign   lane3_r134  =  simd__scntl__lane_r134 [3] ;
  assign   lane3_r135  =  simd__scntl__lane_r135 [3] ;

// Lane 4                 
  assign   lane4_r128  =  simd__scntl__lane_r128 [4] ;
  assign   lane4_r129  =  simd__scntl__lane_r129 [4] ;
  assign   lane4_r130  =  simd__scntl__lane_r130 [4] ;
  assign   lane4_r131  =  simd__scntl__lane_r131 [4] ;
  assign   lane4_r132  =  simd__scntl__lane_r132 [4] ;
  assign   lane4_r133  =  simd__scntl__lane_r133 [4] ;
  assign   lane4_r134  =  simd__scntl__lane_r134 [4] ;
  assign   lane4_r135  =  simd__scntl__lane_r135 [4] ;

// Lane 5                 
  assign   lane5_r128  =  simd__scntl__lane_r128 [5] ;
  assign   lane5_r129  =  simd__scntl__lane_r129 [5] ;
  assign   lane5_r130  =  simd__scntl__lane_r130 [5] ;
  assign   lane5_r131  =  simd__scntl__lane_r131 [5] ;
  assign   lane5_r132  =  simd__scntl__lane_r132 [5] ;
  assign   lane5_r133  =  simd__scntl__lane_r133 [5] ;
  assign   lane5_r134  =  simd__scntl__lane_r134 [5] ;
  assign   lane5_r135  =  simd__scntl__lane_r135 [5] ;

// Lane 6                 
  assign   lane6_r128  =  simd__scntl__lane_r128 [6] ;
  assign   lane6_r129  =  simd__scntl__lane_r129 [6] ;
  assign   lane6_r130  =  simd__scntl__lane_r130 [6] ;
  assign   lane6_r131  =  simd__scntl__lane_r131 [6] ;
  assign   lane6_r132  =  simd__scntl__lane_r132 [6] ;
  assign   lane6_r133  =  simd__scntl__lane_r133 [6] ;
  assign   lane6_r134  =  simd__scntl__lane_r134 [6] ;
  assign   lane6_r135  =  simd__scntl__lane_r135 [6] ;

// Lane 7                 
  assign   lane7_r128  =  simd__scntl__lane_r128 [7] ;
  assign   lane7_r129  =  simd__scntl__lane_r129 [7] ;
  assign   lane7_r130  =  simd__scntl__lane_r130 [7] ;
  assign   lane7_r131  =  simd__scntl__lane_r131 [7] ;
  assign   lane7_r132  =  simd__scntl__lane_r132 [7] ;
  assign   lane7_r133  =  simd__scntl__lane_r133 [7] ;
  assign   lane7_r134  =  simd__scntl__lane_r134 [7] ;
  assign   lane7_r135  =  simd__scntl__lane_r135 [7] ;

// Lane 8                 
  assign   lane8_r128  =  simd__scntl__lane_r128 [8] ;
  assign   lane8_r129  =  simd__scntl__lane_r129 [8] ;
  assign   lane8_r130  =  simd__scntl__lane_r130 [8] ;
  assign   lane8_r131  =  simd__scntl__lane_r131 [8] ;
  assign   lane8_r132  =  simd__scntl__lane_r132 [8] ;
  assign   lane8_r133  =  simd__scntl__lane_r133 [8] ;
  assign   lane8_r134  =  simd__scntl__lane_r134 [8] ;
  assign   lane8_r135  =  simd__scntl__lane_r135 [8] ;

// Lane 9                 
  assign   lane9_r128  =  simd__scntl__lane_r128 [9] ;
  assign   lane9_r129  =  simd__scntl__lane_r129 [9] ;
  assign   lane9_r130  =  simd__scntl__lane_r130 [9] ;
  assign   lane9_r131  =  simd__scntl__lane_r131 [9] ;
  assign   lane9_r132  =  simd__scntl__lane_r132 [9] ;
  assign   lane9_r133  =  simd__scntl__lane_r133 [9] ;
  assign   lane9_r134  =  simd__scntl__lane_r134 [9] ;
  assign   lane9_r135  =  simd__scntl__lane_r135 [9] ;

// Lane 10                 
  assign   lane10_r128  =  simd__scntl__lane_r128 [10] ;
  assign   lane10_r129  =  simd__scntl__lane_r129 [10] ;
  assign   lane10_r130  =  simd__scntl__lane_r130 [10] ;
  assign   lane10_r131  =  simd__scntl__lane_r131 [10] ;
  assign   lane10_r132  =  simd__scntl__lane_r132 [10] ;
  assign   lane10_r133  =  simd__scntl__lane_r133 [10] ;
  assign   lane10_r134  =  simd__scntl__lane_r134 [10] ;
  assign   lane10_r135  =  simd__scntl__lane_r135 [10] ;

// Lane 11                 
  assign   lane11_r128  =  simd__scntl__lane_r128 [11] ;
  assign   lane11_r129  =  simd__scntl__lane_r129 [11] ;
  assign   lane11_r130  =  simd__scntl__lane_r130 [11] ;
  assign   lane11_r131  =  simd__scntl__lane_r131 [11] ;
  assign   lane11_r132  =  simd__scntl__lane_r132 [11] ;
  assign   lane11_r133  =  simd__scntl__lane_r133 [11] ;
  assign   lane11_r134  =  simd__scntl__lane_r134 [11] ;
  assign   lane11_r135  =  simd__scntl__lane_r135 [11] ;

// Lane 12                 
  assign   lane12_r128  =  simd__scntl__lane_r128 [12] ;
  assign   lane12_r129  =  simd__scntl__lane_r129 [12] ;
  assign   lane12_r130  =  simd__scntl__lane_r130 [12] ;
  assign   lane12_r131  =  simd__scntl__lane_r131 [12] ;
  assign   lane12_r132  =  simd__scntl__lane_r132 [12] ;
  assign   lane12_r133  =  simd__scntl__lane_r133 [12] ;
  assign   lane12_r134  =  simd__scntl__lane_r134 [12] ;
  assign   lane12_r135  =  simd__scntl__lane_r135 [12] ;

// Lane 13                 
  assign   lane13_r128  =  simd__scntl__lane_r128 [13] ;
  assign   lane13_r129  =  simd__scntl__lane_r129 [13] ;
  assign   lane13_r130  =  simd__scntl__lane_r130 [13] ;
  assign   lane13_r131  =  simd__scntl__lane_r131 [13] ;
  assign   lane13_r132  =  simd__scntl__lane_r132 [13] ;
  assign   lane13_r133  =  simd__scntl__lane_r133 [13] ;
  assign   lane13_r134  =  simd__scntl__lane_r134 [13] ;
  assign   lane13_r135  =  simd__scntl__lane_r135 [13] ;

// Lane 14                 
  assign   lane14_r128  =  simd__scntl__lane_r128 [14] ;
  assign   lane14_r129  =  simd__scntl__lane_r129 [14] ;
  assign   lane14_r130  =  simd__scntl__lane_r130 [14] ;
  assign   lane14_r131  =  simd__scntl__lane_r131 [14] ;
  assign   lane14_r132  =  simd__scntl__lane_r132 [14] ;
  assign   lane14_r133  =  simd__scntl__lane_r133 [14] ;
  assign   lane14_r134  =  simd__scntl__lane_r134 [14] ;
  assign   lane14_r135  =  simd__scntl__lane_r135 [14] ;

// Lane 15                 
  assign   lane15_r128  =  simd__scntl__lane_r128 [15] ;
  assign   lane15_r129  =  simd__scntl__lane_r129 [15] ;
  assign   lane15_r130  =  simd__scntl__lane_r130 [15] ;
  assign   lane15_r131  =  simd__scntl__lane_r131 [15] ;
  assign   lane15_r132  =  simd__scntl__lane_r132 [15] ;
  assign   lane15_r133  =  simd__scntl__lane_r133 [15] ;
  assign   lane15_r134  =  simd__scntl__lane_r134 [15] ;
  assign   lane15_r135  =  simd__scntl__lane_r135 [15] ;

// Lane 16                 
  assign   lane16_r128  =  simd__scntl__lane_r128 [16] ;
  assign   lane16_r129  =  simd__scntl__lane_r129 [16] ;
  assign   lane16_r130  =  simd__scntl__lane_r130 [16] ;
  assign   lane16_r131  =  simd__scntl__lane_r131 [16] ;
  assign   lane16_r132  =  simd__scntl__lane_r132 [16] ;
  assign   lane16_r133  =  simd__scntl__lane_r133 [16] ;
  assign   lane16_r134  =  simd__scntl__lane_r134 [16] ;
  assign   lane16_r135  =  simd__scntl__lane_r135 [16] ;

// Lane 17                 
  assign   lane17_r128  =  simd__scntl__lane_r128 [17] ;
  assign   lane17_r129  =  simd__scntl__lane_r129 [17] ;
  assign   lane17_r130  =  simd__scntl__lane_r130 [17] ;
  assign   lane17_r131  =  simd__scntl__lane_r131 [17] ;
  assign   lane17_r132  =  simd__scntl__lane_r132 [17] ;
  assign   lane17_r133  =  simd__scntl__lane_r133 [17] ;
  assign   lane17_r134  =  simd__scntl__lane_r134 [17] ;
  assign   lane17_r135  =  simd__scntl__lane_r135 [17] ;

// Lane 18                 
  assign   lane18_r128  =  simd__scntl__lane_r128 [18] ;
  assign   lane18_r129  =  simd__scntl__lane_r129 [18] ;
  assign   lane18_r130  =  simd__scntl__lane_r130 [18] ;
  assign   lane18_r131  =  simd__scntl__lane_r131 [18] ;
  assign   lane18_r132  =  simd__scntl__lane_r132 [18] ;
  assign   lane18_r133  =  simd__scntl__lane_r133 [18] ;
  assign   lane18_r134  =  simd__scntl__lane_r134 [18] ;
  assign   lane18_r135  =  simd__scntl__lane_r135 [18] ;

// Lane 19                 
  assign   lane19_r128  =  simd__scntl__lane_r128 [19] ;
  assign   lane19_r129  =  simd__scntl__lane_r129 [19] ;
  assign   lane19_r130  =  simd__scntl__lane_r130 [19] ;
  assign   lane19_r131  =  simd__scntl__lane_r131 [19] ;
  assign   lane19_r132  =  simd__scntl__lane_r132 [19] ;
  assign   lane19_r133  =  simd__scntl__lane_r133 [19] ;
  assign   lane19_r134  =  simd__scntl__lane_r134 [19] ;
  assign   lane19_r135  =  simd__scntl__lane_r135 [19] ;

// Lane 20                 
  assign   lane20_r128  =  simd__scntl__lane_r128 [20] ;
  assign   lane20_r129  =  simd__scntl__lane_r129 [20] ;
  assign   lane20_r130  =  simd__scntl__lane_r130 [20] ;
  assign   lane20_r131  =  simd__scntl__lane_r131 [20] ;
  assign   lane20_r132  =  simd__scntl__lane_r132 [20] ;
  assign   lane20_r133  =  simd__scntl__lane_r133 [20] ;
  assign   lane20_r134  =  simd__scntl__lane_r134 [20] ;
  assign   lane20_r135  =  simd__scntl__lane_r135 [20] ;

// Lane 21                 
  assign   lane21_r128  =  simd__scntl__lane_r128 [21] ;
  assign   lane21_r129  =  simd__scntl__lane_r129 [21] ;
  assign   lane21_r130  =  simd__scntl__lane_r130 [21] ;
  assign   lane21_r131  =  simd__scntl__lane_r131 [21] ;
  assign   lane21_r132  =  simd__scntl__lane_r132 [21] ;
  assign   lane21_r133  =  simd__scntl__lane_r133 [21] ;
  assign   lane21_r134  =  simd__scntl__lane_r134 [21] ;
  assign   lane21_r135  =  simd__scntl__lane_r135 [21] ;

// Lane 22                 
  assign   lane22_r128  =  simd__scntl__lane_r128 [22] ;
  assign   lane22_r129  =  simd__scntl__lane_r129 [22] ;
  assign   lane22_r130  =  simd__scntl__lane_r130 [22] ;
  assign   lane22_r131  =  simd__scntl__lane_r131 [22] ;
  assign   lane22_r132  =  simd__scntl__lane_r132 [22] ;
  assign   lane22_r133  =  simd__scntl__lane_r133 [22] ;
  assign   lane22_r134  =  simd__scntl__lane_r134 [22] ;
  assign   lane22_r135  =  simd__scntl__lane_r135 [22] ;

// Lane 23                 
  assign   lane23_r128  =  simd__scntl__lane_r128 [23] ;
  assign   lane23_r129  =  simd__scntl__lane_r129 [23] ;
  assign   lane23_r130  =  simd__scntl__lane_r130 [23] ;
  assign   lane23_r131  =  simd__scntl__lane_r131 [23] ;
  assign   lane23_r132  =  simd__scntl__lane_r132 [23] ;
  assign   lane23_r133  =  simd__scntl__lane_r133 [23] ;
  assign   lane23_r134  =  simd__scntl__lane_r134 [23] ;
  assign   lane23_r135  =  simd__scntl__lane_r135 [23] ;

// Lane 24                 
  assign   lane24_r128  =  simd__scntl__lane_r128 [24] ;
  assign   lane24_r129  =  simd__scntl__lane_r129 [24] ;
  assign   lane24_r130  =  simd__scntl__lane_r130 [24] ;
  assign   lane24_r131  =  simd__scntl__lane_r131 [24] ;
  assign   lane24_r132  =  simd__scntl__lane_r132 [24] ;
  assign   lane24_r133  =  simd__scntl__lane_r133 [24] ;
  assign   lane24_r134  =  simd__scntl__lane_r134 [24] ;
  assign   lane24_r135  =  simd__scntl__lane_r135 [24] ;

// Lane 25                 
  assign   lane25_r128  =  simd__scntl__lane_r128 [25] ;
  assign   lane25_r129  =  simd__scntl__lane_r129 [25] ;
  assign   lane25_r130  =  simd__scntl__lane_r130 [25] ;
  assign   lane25_r131  =  simd__scntl__lane_r131 [25] ;
  assign   lane25_r132  =  simd__scntl__lane_r132 [25] ;
  assign   lane25_r133  =  simd__scntl__lane_r133 [25] ;
  assign   lane25_r134  =  simd__scntl__lane_r134 [25] ;
  assign   lane25_r135  =  simd__scntl__lane_r135 [25] ;

// Lane 26                 
  assign   lane26_r128  =  simd__scntl__lane_r128 [26] ;
  assign   lane26_r129  =  simd__scntl__lane_r129 [26] ;
  assign   lane26_r130  =  simd__scntl__lane_r130 [26] ;
  assign   lane26_r131  =  simd__scntl__lane_r131 [26] ;
  assign   lane26_r132  =  simd__scntl__lane_r132 [26] ;
  assign   lane26_r133  =  simd__scntl__lane_r133 [26] ;
  assign   lane26_r134  =  simd__scntl__lane_r134 [26] ;
  assign   lane26_r135  =  simd__scntl__lane_r135 [26] ;

// Lane 27                 
  assign   lane27_r128  =  simd__scntl__lane_r128 [27] ;
  assign   lane27_r129  =  simd__scntl__lane_r129 [27] ;
  assign   lane27_r130  =  simd__scntl__lane_r130 [27] ;
  assign   lane27_r131  =  simd__scntl__lane_r131 [27] ;
  assign   lane27_r132  =  simd__scntl__lane_r132 [27] ;
  assign   lane27_r133  =  simd__scntl__lane_r133 [27] ;
  assign   lane27_r134  =  simd__scntl__lane_r134 [27] ;
  assign   lane27_r135  =  simd__scntl__lane_r135 [27] ;

// Lane 28                 
  assign   lane28_r128  =  simd__scntl__lane_r128 [28] ;
  assign   lane28_r129  =  simd__scntl__lane_r129 [28] ;
  assign   lane28_r130  =  simd__scntl__lane_r130 [28] ;
  assign   lane28_r131  =  simd__scntl__lane_r131 [28] ;
  assign   lane28_r132  =  simd__scntl__lane_r132 [28] ;
  assign   lane28_r133  =  simd__scntl__lane_r133 [28] ;
  assign   lane28_r134  =  simd__scntl__lane_r134 [28] ;
  assign   lane28_r135  =  simd__scntl__lane_r135 [28] ;

// Lane 29                 
  assign   lane29_r128  =  simd__scntl__lane_r128 [29] ;
  assign   lane29_r129  =  simd__scntl__lane_r129 [29] ;
  assign   lane29_r130  =  simd__scntl__lane_r130 [29] ;
  assign   lane29_r131  =  simd__scntl__lane_r131 [29] ;
  assign   lane29_r132  =  simd__scntl__lane_r132 [29] ;
  assign   lane29_r133  =  simd__scntl__lane_r133 [29] ;
  assign   lane29_r134  =  simd__scntl__lane_r134 [29] ;
  assign   lane29_r135  =  simd__scntl__lane_r135 [29] ;

// Lane 30                 
  assign   lane30_r128  =  simd__scntl__lane_r128 [30] ;
  assign   lane30_r129  =  simd__scntl__lane_r129 [30] ;
  assign   lane30_r130  =  simd__scntl__lane_r130 [30] ;
  assign   lane30_r131  =  simd__scntl__lane_r131 [30] ;
  assign   lane30_r132  =  simd__scntl__lane_r132 [30] ;
  assign   lane30_r133  =  simd__scntl__lane_r133 [30] ;
  assign   lane30_r134  =  simd__scntl__lane_r134 [30] ;
  assign   lane30_r135  =  simd__scntl__lane_r135 [30] ;

// Lane 31                 
  assign   lane31_r128  =  simd__scntl__lane_r128 [31] ;
  assign   lane31_r129  =  simd__scntl__lane_r129 [31] ;
  assign   lane31_r130  =  simd__scntl__lane_r130 [31] ;
  assign   lane31_r131  =  simd__scntl__lane_r131 [31] ;
  assign   lane31_r132  =  simd__scntl__lane_r132 [31] ;
  assign   lane31_r133  =  simd__scntl__lane_r133 [31] ;
  assign   lane31_r134  =  simd__scntl__lane_r134 [31] ;
  assign   lane31_r135  =  simd__scntl__lane_r135 [31] ;
