
    output                                         stu__mgr0__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr0__cntl           ;
    input                                          mgr0__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr0__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr0__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr0__oob_data       ;

    input                                          pe0__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe0__stu__cntl           ;
    output                                         stu__pe0__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe0__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe0__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe0__stu__oob_data       ;

    output                                         stu__mgr1__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr1__cntl           ;
    input                                          mgr1__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr1__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr1__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr1__oob_data       ;

    input                                          pe1__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe1__stu__cntl           ;
    output                                         stu__pe1__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe1__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe1__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe1__stu__oob_data       ;

    output                                         stu__mgr2__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr2__cntl           ;
    input                                          mgr2__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr2__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr2__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr2__oob_data       ;

    input                                          pe2__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe2__stu__cntl           ;
    output                                         stu__pe2__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe2__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe2__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe2__stu__oob_data       ;

    output                                         stu__mgr3__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr3__cntl           ;
    input                                          mgr3__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr3__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr3__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr3__oob_data       ;

    input                                          pe3__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe3__stu__cntl           ;
    output                                         stu__pe3__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe3__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe3__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe3__stu__oob_data       ;

