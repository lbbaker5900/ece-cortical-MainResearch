
   reg [`PE_PE_ID_BITMASK_RANGE      ] thisPeBitMask       ; 