

            // DMA port 0
            dma__memc__write_valid0 ,
            dma__memc__write_address0 ,
            dma__memc__write_data0 ,
            memc__dma__write_ready0 ,
            dma__memc__read_valid0 ,
            dma__memc__read_address0 ,
            memc__dma__read_data0 ,
            memc__dma__read_data_valid0 ,
            memc__dma__read_ready0 ,
            dma__memc__read_pause0 ,

            // DMA port 1
            dma__memc__write_valid1 ,
            dma__memc__write_address1 ,
            dma__memc__write_data1 ,
            memc__dma__write_ready1 ,
            dma__memc__read_valid1 ,
            dma__memc__read_address1 ,
            memc__dma__read_data1 ,
            memc__dma__read_data_valid1 ,
            memc__dma__read_ready1 ,
            dma__memc__read_pause1 ,

            // DMA port 2
            dma__memc__write_valid2 ,
            dma__memc__write_address2 ,
            dma__memc__write_data2 ,
            memc__dma__write_ready2 ,
            dma__memc__read_valid2 ,
            dma__memc__read_address2 ,
            memc__dma__read_data2 ,
            memc__dma__read_data_valid2 ,
            memc__dma__read_ready2 ,
            dma__memc__read_pause2 ,

            // DMA port 3
            dma__memc__write_valid3 ,
            dma__memc__write_address3 ,
            dma__memc__write_data3 ,
            memc__dma__write_ready3 ,
            dma__memc__read_valid3 ,
            dma__memc__read_address3 ,
            memc__dma__read_data3 ,
            memc__dma__read_data_valid3 ,
            memc__dma__read_ready3 ,
            dma__memc__read_pause3 ,

            // DMA port 4
            dma__memc__write_valid4 ,
            dma__memc__write_address4 ,
            dma__memc__write_data4 ,
            memc__dma__write_ready4 ,
            dma__memc__read_valid4 ,
            dma__memc__read_address4 ,
            memc__dma__read_data4 ,
            memc__dma__read_data_valid4 ,
            memc__dma__read_ready4 ,
            dma__memc__read_pause4 ,

            // DMA port 5
            dma__memc__write_valid5 ,
            dma__memc__write_address5 ,
            dma__memc__write_data5 ,
            memc__dma__write_ready5 ,
            dma__memc__read_valid5 ,
            dma__memc__read_address5 ,
            memc__dma__read_data5 ,
            memc__dma__read_data_valid5 ,
            memc__dma__read_ready5 ,
            dma__memc__read_pause5 ,

            // DMA port 6
            dma__memc__write_valid6 ,
            dma__memc__write_address6 ,
            dma__memc__write_data6 ,
            memc__dma__write_ready6 ,
            dma__memc__read_valid6 ,
            dma__memc__read_address6 ,
            memc__dma__read_data6 ,
            memc__dma__read_data_valid6 ,
            memc__dma__read_ready6 ,
            dma__memc__read_pause6 ,

            // DMA port 7
            dma__memc__write_valid7 ,
            dma__memc__write_address7 ,
            dma__memc__write_data7 ,
            memc__dma__write_ready7 ,
            dma__memc__read_valid7 ,
            dma__memc__read_address7 ,
            memc__dma__read_data7 ,
            memc__dma__read_data_valid7 ,
            memc__dma__read_ready7 ,
            dma__memc__read_pause7 ,

            // DMA port 8
            dma__memc__write_valid8 ,
            dma__memc__write_address8 ,
            dma__memc__write_data8 ,
            memc__dma__write_ready8 ,
            dma__memc__read_valid8 ,
            dma__memc__read_address8 ,
            memc__dma__read_data8 ,
            memc__dma__read_data_valid8 ,
            memc__dma__read_ready8 ,
            dma__memc__read_pause8 ,

            // DMA port 9
            dma__memc__write_valid9 ,
            dma__memc__write_address9 ,
            dma__memc__write_data9 ,
            memc__dma__write_ready9 ,
            dma__memc__read_valid9 ,
            dma__memc__read_address9 ,
            memc__dma__read_data9 ,
            memc__dma__read_data_valid9 ,
            memc__dma__read_ready9 ,
            dma__memc__read_pause9 ,

            // DMA port 10
            dma__memc__write_valid10 ,
            dma__memc__write_address10 ,
            dma__memc__write_data10 ,
            memc__dma__write_ready10 ,
            dma__memc__read_valid10 ,
            dma__memc__read_address10 ,
            memc__dma__read_data10 ,
            memc__dma__read_data_valid10 ,
            memc__dma__read_ready10 ,
            dma__memc__read_pause10 ,

            // DMA port 11
            dma__memc__write_valid11 ,
            dma__memc__write_address11 ,
            dma__memc__write_data11 ,
            memc__dma__write_ready11 ,
            dma__memc__read_valid11 ,
            dma__memc__read_address11 ,
            memc__dma__read_data11 ,
            memc__dma__read_data_valid11 ,
            memc__dma__read_ready11 ,
            dma__memc__read_pause11 ,

            // DMA port 12
            dma__memc__write_valid12 ,
            dma__memc__write_address12 ,
            dma__memc__write_data12 ,
            memc__dma__write_ready12 ,
            dma__memc__read_valid12 ,
            dma__memc__read_address12 ,
            memc__dma__read_data12 ,
            memc__dma__read_data_valid12 ,
            memc__dma__read_ready12 ,
            dma__memc__read_pause12 ,

            // DMA port 13
            dma__memc__write_valid13 ,
            dma__memc__write_address13 ,
            dma__memc__write_data13 ,
            memc__dma__write_ready13 ,
            dma__memc__read_valid13 ,
            dma__memc__read_address13 ,
            memc__dma__read_data13 ,
            memc__dma__read_data_valid13 ,
            memc__dma__read_ready13 ,
            dma__memc__read_pause13 ,

            // DMA port 14
            dma__memc__write_valid14 ,
            dma__memc__write_address14 ,
            dma__memc__write_data14 ,
            memc__dma__write_ready14 ,
            dma__memc__read_valid14 ,
            dma__memc__read_address14 ,
            memc__dma__read_data14 ,
            memc__dma__read_data_valid14 ,
            memc__dma__read_ready14 ,
            dma__memc__read_pause14 ,

            // DMA port 15
            dma__memc__write_valid15 ,
            dma__memc__write_address15 ,
            dma__memc__write_data15 ,
            memc__dma__write_ready15 ,
            dma__memc__read_valid15 ,
            dma__memc__read_address15 ,
            memc__dma__read_data15 ,
            memc__dma__read_data_valid15 ,
            memc__dma__read_ready15 ,
            dma__memc__read_pause15 ,

            // DMA port 16
            dma__memc__write_valid16 ,
            dma__memc__write_address16 ,
            dma__memc__write_data16 ,
            memc__dma__write_ready16 ,
            dma__memc__read_valid16 ,
            dma__memc__read_address16 ,
            memc__dma__read_data16 ,
            memc__dma__read_data_valid16 ,
            memc__dma__read_ready16 ,
            dma__memc__read_pause16 ,

            // DMA port 17
            dma__memc__write_valid17 ,
            dma__memc__write_address17 ,
            dma__memc__write_data17 ,
            memc__dma__write_ready17 ,
            dma__memc__read_valid17 ,
            dma__memc__read_address17 ,
            memc__dma__read_data17 ,
            memc__dma__read_data_valid17 ,
            memc__dma__read_ready17 ,
            dma__memc__read_pause17 ,

            // DMA port 18
            dma__memc__write_valid18 ,
            dma__memc__write_address18 ,
            dma__memc__write_data18 ,
            memc__dma__write_ready18 ,
            dma__memc__read_valid18 ,
            dma__memc__read_address18 ,
            memc__dma__read_data18 ,
            memc__dma__read_data_valid18 ,
            memc__dma__read_ready18 ,
            dma__memc__read_pause18 ,

            // DMA port 19
            dma__memc__write_valid19 ,
            dma__memc__write_address19 ,
            dma__memc__write_data19 ,
            memc__dma__write_ready19 ,
            dma__memc__read_valid19 ,
            dma__memc__read_address19 ,
            memc__dma__read_data19 ,
            memc__dma__read_data_valid19 ,
            memc__dma__read_ready19 ,
            dma__memc__read_pause19 ,

            // DMA port 20
            dma__memc__write_valid20 ,
            dma__memc__write_address20 ,
            dma__memc__write_data20 ,
            memc__dma__write_ready20 ,
            dma__memc__read_valid20 ,
            dma__memc__read_address20 ,
            memc__dma__read_data20 ,
            memc__dma__read_data_valid20 ,
            memc__dma__read_ready20 ,
            dma__memc__read_pause20 ,

            // DMA port 21
            dma__memc__write_valid21 ,
            dma__memc__write_address21 ,
            dma__memc__write_data21 ,
            memc__dma__write_ready21 ,
            dma__memc__read_valid21 ,
            dma__memc__read_address21 ,
            memc__dma__read_data21 ,
            memc__dma__read_data_valid21 ,
            memc__dma__read_ready21 ,
            dma__memc__read_pause21 ,

            // DMA port 22
            dma__memc__write_valid22 ,
            dma__memc__write_address22 ,
            dma__memc__write_data22 ,
            memc__dma__write_ready22 ,
            dma__memc__read_valid22 ,
            dma__memc__read_address22 ,
            memc__dma__read_data22 ,
            memc__dma__read_data_valid22 ,
            memc__dma__read_ready22 ,
            dma__memc__read_pause22 ,

            // DMA port 23
            dma__memc__write_valid23 ,
            dma__memc__write_address23 ,
            dma__memc__write_data23 ,
            memc__dma__write_ready23 ,
            dma__memc__read_valid23 ,
            dma__memc__read_address23 ,
            memc__dma__read_data23 ,
            memc__dma__read_data_valid23 ,
            memc__dma__read_ready23 ,
            dma__memc__read_pause23 ,

            // DMA port 24
            dma__memc__write_valid24 ,
            dma__memc__write_address24 ,
            dma__memc__write_data24 ,
            memc__dma__write_ready24 ,
            dma__memc__read_valid24 ,
            dma__memc__read_address24 ,
            memc__dma__read_data24 ,
            memc__dma__read_data_valid24 ,
            memc__dma__read_ready24 ,
            dma__memc__read_pause24 ,

            // DMA port 25
            dma__memc__write_valid25 ,
            dma__memc__write_address25 ,
            dma__memc__write_data25 ,
            memc__dma__write_ready25 ,
            dma__memc__read_valid25 ,
            dma__memc__read_address25 ,
            memc__dma__read_data25 ,
            memc__dma__read_data_valid25 ,
            memc__dma__read_ready25 ,
            dma__memc__read_pause25 ,

            // DMA port 26
            dma__memc__write_valid26 ,
            dma__memc__write_address26 ,
            dma__memc__write_data26 ,
            memc__dma__write_ready26 ,
            dma__memc__read_valid26 ,
            dma__memc__read_address26 ,
            memc__dma__read_data26 ,
            memc__dma__read_data_valid26 ,
            memc__dma__read_ready26 ,
            dma__memc__read_pause26 ,

            // DMA port 27
            dma__memc__write_valid27 ,
            dma__memc__write_address27 ,
            dma__memc__write_data27 ,
            memc__dma__write_ready27 ,
            dma__memc__read_valid27 ,
            dma__memc__read_address27 ,
            memc__dma__read_data27 ,
            memc__dma__read_data_valid27 ,
            memc__dma__read_ready27 ,
            dma__memc__read_pause27 ,

            // DMA port 28
            dma__memc__write_valid28 ,
            dma__memc__write_address28 ,
            dma__memc__write_data28 ,
            memc__dma__write_ready28 ,
            dma__memc__read_valid28 ,
            dma__memc__read_address28 ,
            memc__dma__read_data28 ,
            memc__dma__read_data_valid28 ,
            memc__dma__read_ready28 ,
            dma__memc__read_pause28 ,

            // DMA port 29
            dma__memc__write_valid29 ,
            dma__memc__write_address29 ,
            dma__memc__write_data29 ,
            memc__dma__write_ready29 ,
            dma__memc__read_valid29 ,
            dma__memc__read_address29 ,
            memc__dma__read_data29 ,
            memc__dma__read_data_valid29 ,
            memc__dma__read_ready29 ,
            dma__memc__read_pause29 ,

            // DMA port 30
            dma__memc__write_valid30 ,
            dma__memc__write_address30 ,
            dma__memc__write_data30 ,
            memc__dma__write_ready30 ,
            dma__memc__read_valid30 ,
            dma__memc__read_address30 ,
            memc__dma__read_data30 ,
            memc__dma__read_data_valid30 ,
            memc__dma__read_ready30 ,
            dma__memc__read_pause30 ,

            // DMA port 31
            dma__memc__write_valid31 ,
            dma__memc__write_address31 ,
            dma__memc__write_data31 ,
            memc__dma__write_ready31 ,
            dma__memc__read_valid31 ,
            dma__memc__read_address31 ,
            memc__dma__read_data31 ,
            memc__dma__read_data_valid31 ,
            memc__dma__read_ready31 ,
            dma__memc__read_pause31 ,
