

            // ##################################################
            // Memory Stream Source addresses

            // Stream 0 Source address
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [0] = 32'b000000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [1] = 32'b000000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [2] = 32'b000000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [3] = 32'b000000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [4] = 32'b000000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [5] = 32'b000000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [6] = 32'b000000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [7] = 32'b000000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [8] = 32'b000000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [9] = 32'b000000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [10] = 32'b000000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [11] = 32'b000000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [12] = 32'b000000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [13] = 32'b000000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [14] = 32'b000000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [15] = 32'b000000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [16] = 32'b000000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [17] = 32'b000000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [18] = 32'b000000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [19] = 32'b000000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [20] = 32'b000000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [21] = 32'b000000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [22] = 32'b000000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [23] = 32'b000000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [24] = 32'b000000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [25] = 32'b000000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [26] = 32'b000000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [27] = 32'b000000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [28] = 32'b000000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [29] = 32'b000000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [30] = 32'b000000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [31] = 32'b000000_11111__0_0000_1000_0000;
            // Stream 1 Source address
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [0] = 32'b000000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [1] = 32'b000000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [2] = 32'b000000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [3] = 32'b000000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [4] = 32'b000000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [5] = 32'b000000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [6] = 32'b000000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [7] = 32'b000000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [8] = 32'b000000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [9] = 32'b000000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [10] = 32'b000000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [11] = 32'b000000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [12] = 32'b000000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [13] = 32'b000000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [14] = 32'b000000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [15] = 32'b000000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [16] = 32'b000000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [17] = 32'b000000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [18] = 32'b000000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [19] = 32'b000000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [20] = 32'b000000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [21] = 32'b000000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [22] = 32'b000000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [23] = 32'b000000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [24] = 32'b000000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [25] = 32'b000000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [26] = 32'b000000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [27] = 32'b000000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [28] = 32'b000000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [29] = 32'b000000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [30] = 32'b000000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [31] = 32'b000000_11111__0_1000_0000_0000;
            // Stream 0 Source address
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [0] = 32'b000001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [1] = 32'b000001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [2] = 32'b000001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [3] = 32'b000001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [4] = 32'b000001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [5] = 32'b000001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [6] = 32'b000001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [7] = 32'b000001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [8] = 32'b000001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [9] = 32'b000001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [10] = 32'b000001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [11] = 32'b000001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [12] = 32'b000001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [13] = 32'b000001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [14] = 32'b000001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [15] = 32'b000001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [16] = 32'b000001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [17] = 32'b000001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [18] = 32'b000001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [19] = 32'b000001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [20] = 32'b000001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [21] = 32'b000001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [22] = 32'b000001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [23] = 32'b000001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [24] = 32'b000001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [25] = 32'b000001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [26] = 32'b000001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [27] = 32'b000001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [28] = 32'b000001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [29] = 32'b000001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [30] = 32'b000001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [31] = 32'b000001_11111__0_0000_1000_0000;
            // Stream 1 Source address
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [0] = 32'b000001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [1] = 32'b000001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [2] = 32'b000001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [3] = 32'b000001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [4] = 32'b000001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [5] = 32'b000001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [6] = 32'b000001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [7] = 32'b000001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [8] = 32'b000001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [9] = 32'b000001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [10] = 32'b000001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [11] = 32'b000001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [12] = 32'b000001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [13] = 32'b000001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [14] = 32'b000001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [15] = 32'b000001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [16] = 32'b000001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [17] = 32'b000001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [18] = 32'b000001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [19] = 32'b000001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [20] = 32'b000001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [21] = 32'b000001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [22] = 32'b000001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [23] = 32'b000001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [24] = 32'b000001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [25] = 32'b000001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [26] = 32'b000001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [27] = 32'b000001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [28] = 32'b000001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [29] = 32'b000001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [30] = 32'b000001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [31] = 32'b000001_11111__0_1000_0000_0000;
            // Stream 0 Source address
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [0] = 32'b000010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [1] = 32'b000010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [2] = 32'b000010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [3] = 32'b000010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [4] = 32'b000010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [5] = 32'b000010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [6] = 32'b000010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [7] = 32'b000010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [8] = 32'b000010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [9] = 32'b000010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [10] = 32'b000010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [11] = 32'b000010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [12] = 32'b000010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [13] = 32'b000010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [14] = 32'b000010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [15] = 32'b000010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [16] = 32'b000010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [17] = 32'b000010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [18] = 32'b000010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [19] = 32'b000010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [20] = 32'b000010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [21] = 32'b000010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [22] = 32'b000010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [23] = 32'b000010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [24] = 32'b000010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [25] = 32'b000010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [26] = 32'b000010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [27] = 32'b000010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [28] = 32'b000010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [29] = 32'b000010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [30] = 32'b000010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [31] = 32'b000010_11111__0_0000_1000_0000;
            // Stream 1 Source address
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [0] = 32'b000010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [1] = 32'b000010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [2] = 32'b000010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [3] = 32'b000010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [4] = 32'b000010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [5] = 32'b000010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [6] = 32'b000010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [7] = 32'b000010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [8] = 32'b000010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [9] = 32'b000010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [10] = 32'b000010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [11] = 32'b000010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [12] = 32'b000010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [13] = 32'b000010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [14] = 32'b000010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [15] = 32'b000010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [16] = 32'b000010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [17] = 32'b000010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [18] = 32'b000010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [19] = 32'b000010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [20] = 32'b000010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [21] = 32'b000010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [22] = 32'b000010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [23] = 32'b000010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [24] = 32'b000010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [25] = 32'b000010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [26] = 32'b000010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [27] = 32'b000010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [28] = 32'b000010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [29] = 32'b000010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [30] = 32'b000010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [31] = 32'b000010_11111__0_1000_0000_0000;
            // Stream 0 Source address
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [0] = 32'b000011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [1] = 32'b000011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [2] = 32'b000011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [3] = 32'b000011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [4] = 32'b000011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [5] = 32'b000011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [6] = 32'b000011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [7] = 32'b000011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [8] = 32'b000011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [9] = 32'b000011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [10] = 32'b000011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [11] = 32'b000011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [12] = 32'b000011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [13] = 32'b000011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [14] = 32'b000011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [15] = 32'b000011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [16] = 32'b000011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [17] = 32'b000011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [18] = 32'b000011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [19] = 32'b000011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [20] = 32'b000011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [21] = 32'b000011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [22] = 32'b000011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [23] = 32'b000011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [24] = 32'b000011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [25] = 32'b000011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [26] = 32'b000011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [27] = 32'b000011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [28] = 32'b000011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [29] = 32'b000011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [30] = 32'b000011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [31] = 32'b000011_11111__0_0000_1000_0000;
            // Stream 1 Source address
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [0] = 32'b000011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [1] = 32'b000011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [2] = 32'b000011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [3] = 32'b000011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [4] = 32'b000011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [5] = 32'b000011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [6] = 32'b000011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [7] = 32'b000011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [8] = 32'b000011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [9] = 32'b000011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [10] = 32'b000011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [11] = 32'b000011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [12] = 32'b000011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [13] = 32'b000011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [14] = 32'b000011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [15] = 32'b000011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [16] = 32'b000011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [17] = 32'b000011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [18] = 32'b000011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [19] = 32'b000011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [20] = 32'b000011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [21] = 32'b000011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [22] = 32'b000011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [23] = 32'b000011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [24] = 32'b000011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [25] = 32'b000011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [26] = 32'b000011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [27] = 32'b000011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [28] = 32'b000011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [29] = 32'b000011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [30] = 32'b000011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [31] = 32'b000011_11111__0_1000_0000_0000;


            // ##################################################
            // Memory Destination addresses

            // Stream 0 Destination address
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [0] = 32'b000000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [1] = 32'b000000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [2] = 32'b000000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [3] = 32'b000000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [4] = 32'b000000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [5] = 32'b000000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [6] = 32'b000000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [7] = 32'b000000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [8] = 32'b000000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [9] = 32'b000000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [10] = 32'b000000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [11] = 32'b000000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [12] = 32'b000000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [13] = 32'b000000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [14] = 32'b000000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [15] = 32'b000000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [16] = 32'b000000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [17] = 32'b000000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [18] = 32'b000000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [19] = 32'b000000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [20] = 32'b000000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [21] = 32'b000000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [22] = 32'b000000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [23] = 32'b000000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [24] = 32'b000000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [25] = 32'b000000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [26] = 32'b000000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [27] = 32'b000000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [28] = 32'b000000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [29] = 32'b000000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [30] = 32'b000000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [31] = 32'b000000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [0] = 32'b000000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [1] = 32'b000000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [2] = 32'b000000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [3] = 32'b000000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [4] = 32'b000000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [5] = 32'b000000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [6] = 32'b000000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [7] = 32'b000000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [8] = 32'b000000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [9] = 32'b000000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [10] = 32'b000000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [11] = 32'b000000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [12] = 32'b000000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [13] = 32'b000000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [14] = 32'b000000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [15] = 32'b000000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [16] = 32'b000000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [17] = 32'b000000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [18] = 32'b000000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [19] = 32'b000000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [20] = 32'b000000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [21] = 32'b000000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [22] = 32'b000000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [23] = 32'b000000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [24] = 32'b000000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [25] = 32'b000000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [26] = 32'b000000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [27] = 32'b000000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [28] = 32'b000000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [29] = 32'b000000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [30] = 32'b000000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [31] = 32'b000000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [0] = 32'b000001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [1] = 32'b000001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [2] = 32'b000001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [3] = 32'b000001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [4] = 32'b000001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [5] = 32'b000001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [6] = 32'b000001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [7] = 32'b000001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [8] = 32'b000001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [9] = 32'b000001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [10] = 32'b000001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [11] = 32'b000001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [12] = 32'b000001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [13] = 32'b000001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [14] = 32'b000001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [15] = 32'b000001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [16] = 32'b000001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [17] = 32'b000001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [18] = 32'b000001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [19] = 32'b000001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [20] = 32'b000001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [21] = 32'b000001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [22] = 32'b000001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [23] = 32'b000001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [24] = 32'b000001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [25] = 32'b000001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [26] = 32'b000001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [27] = 32'b000001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [28] = 32'b000001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [29] = 32'b000001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [30] = 32'b000001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [31] = 32'b000001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [0] = 32'b000001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [1] = 32'b000001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [2] = 32'b000001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [3] = 32'b000001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [4] = 32'b000001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [5] = 32'b000001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [6] = 32'b000001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [7] = 32'b000001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [8] = 32'b000001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [9] = 32'b000001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [10] = 32'b000001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [11] = 32'b000001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [12] = 32'b000001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [13] = 32'b000001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [14] = 32'b000001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [15] = 32'b000001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [16] = 32'b000001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [17] = 32'b000001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [18] = 32'b000001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [19] = 32'b000001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [20] = 32'b000001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [21] = 32'b000001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [22] = 32'b000001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [23] = 32'b000001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [24] = 32'b000001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [25] = 32'b000001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [26] = 32'b000001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [27] = 32'b000001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [28] = 32'b000001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [29] = 32'b000001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [30] = 32'b000001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [31] = 32'b000001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [0] = 32'b000010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [1] = 32'b000010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [2] = 32'b000010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [3] = 32'b000010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [4] = 32'b000010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [5] = 32'b000010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [6] = 32'b000010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [7] = 32'b000010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [8] = 32'b000010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [9] = 32'b000010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [10] = 32'b000010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [11] = 32'b000010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [12] = 32'b000010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [13] = 32'b000010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [14] = 32'b000010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [15] = 32'b000010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [16] = 32'b000010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [17] = 32'b000010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [18] = 32'b000010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [19] = 32'b000010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [20] = 32'b000010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [21] = 32'b000010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [22] = 32'b000010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [23] = 32'b000010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [24] = 32'b000010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [25] = 32'b000010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [26] = 32'b000010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [27] = 32'b000010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [28] = 32'b000010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [29] = 32'b000010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [30] = 32'b000010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [31] = 32'b000010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [0] = 32'b000010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [1] = 32'b000010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [2] = 32'b000010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [3] = 32'b000010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [4] = 32'b000010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [5] = 32'b000010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [6] = 32'b000010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [7] = 32'b000010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [8] = 32'b000010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [9] = 32'b000010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [10] = 32'b000010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [11] = 32'b000010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [12] = 32'b000010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [13] = 32'b000010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [14] = 32'b000010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [15] = 32'b000010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [16] = 32'b000010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [17] = 32'b000010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [18] = 32'b000010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [19] = 32'b000010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [20] = 32'b000010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [21] = 32'b000010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [22] = 32'b000010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [23] = 32'b000010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [24] = 32'b000010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [25] = 32'b000010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [26] = 32'b000010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [27] = 32'b000010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [28] = 32'b000010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [29] = 32'b000010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [30] = 32'b000010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [31] = 32'b000010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [0] = 32'b000011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [1] = 32'b000011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [2] = 32'b000011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [3] = 32'b000011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [4] = 32'b000011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [5] = 32'b000011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [6] = 32'b000011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [7] = 32'b000011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [8] = 32'b000011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [9] = 32'b000011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [10] = 32'b000011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [11] = 32'b000011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [12] = 32'b000011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [13] = 32'b000011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [14] = 32'b000011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [15] = 32'b000011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [16] = 32'b000011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [17] = 32'b000011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [18] = 32'b000011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [19] = 32'b000011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [20] = 32'b000011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [21] = 32'b000011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [22] = 32'b000011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [23] = 32'b000011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [24] = 32'b000011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [25] = 32'b000011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [26] = 32'b000011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [27] = 32'b000011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [28] = 32'b000011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [29] = 32'b000011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [30] = 32'b000011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [31] = 32'b000011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [0] = 32'b000011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [1] = 32'b000011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [2] = 32'b000011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [3] = 32'b000011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [4] = 32'b000011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [5] = 32'b000011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [6] = 32'b000011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [7] = 32'b000011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [8] = 32'b000011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [9] = 32'b000011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [10] = 32'b000011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [11] = 32'b000011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [12] = 32'b000011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [13] = 32'b000011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [14] = 32'b000011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [15] = 32'b000011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [16] = 32'b000011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [17] = 32'b000011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [18] = 32'b000011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [19] = 32'b000011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [20] = 32'b000011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [21] = 32'b000011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [22] = 32'b000011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [23] = 32'b000011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [24] = 32'b000011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [25] = 32'b000011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [26] = 32'b000011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [27] = 32'b000011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [28] = 32'b000011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [29] = 32'b000011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [30] = 32'b000011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [31] = 32'b000011_11111__0_1000_0000_0000;

            // ##################################################
            // DMA Type and length of stream

            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;


            // ##################################################
            // Enable and set transfer type

            repeat(10) @(negedge clk); 

            // Enable
            force pe_array_inst.pe_inst[0].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[1].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[2].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[3].pe.rs0[0]           = 1'b1;

            // Operation
            force pe_array_inst.pe_inst[0].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_MEM_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[1].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_MEM_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[2].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_MEM_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[3].pe.rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_MEM_STD_FP_MAC_TO_MEM ;

            repeat(50) @(negedge clk);