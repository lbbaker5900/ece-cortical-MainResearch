`ifndef _wu_fetch_vh
`define _wu_fetch_vh

/*****************************************************************

    File name   : wu_fetch.vh
    Author      : Lee Baker
    Affiliation : North Carolina State University, Raleigh, NC
    Date        : Mar 2017
    email       : lbbaker@ncsu.edu

*****************************************************************/



`endif
