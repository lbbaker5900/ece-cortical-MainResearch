
    output                                         pe0__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe0__stu__cntl           ;
    input                                          stu__pe0__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe0__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe0__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe0__stu__oob_data       ;

    output                                         pe1__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe1__stu__cntl           ;
    input                                          stu__pe1__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe1__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe1__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe1__stu__oob_data       ;

    output                                         pe2__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe2__stu__cntl           ;
    input                                          stu__pe2__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe2__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe2__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe2__stu__oob_data       ;

    output                                         pe3__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe3__stu__cntl           ;
    input                                          stu__pe3__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe3__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe3__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe3__stu__oob_data       ;

