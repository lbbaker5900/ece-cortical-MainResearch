
            // General control and status                  
            .sys__pe0__allSynchronized                  ( sys__pe0__allSynchronized   ),
            .pe0__sys__thisSynchronized                 ( pe0__sys__thisSynchronized  ),
            .pe0__sys__ready                            ( pe0__sys__ready             ),
            .pe0__sys__complete                         ( pe0__sys__complete          ),
            // General control and status                  
            .sys__pe1__allSynchronized                  ( sys__pe1__allSynchronized   ),
            .pe1__sys__thisSynchronized                 ( pe1__sys__thisSynchronized  ),
            .pe1__sys__ready                            ( pe1__sys__ready             ),
            .pe1__sys__complete                         ( pe1__sys__complete          ),
            // General control and status                  
            .sys__pe2__allSynchronized                  ( sys__pe2__allSynchronized   ),
            .pe2__sys__thisSynchronized                 ( pe2__sys__thisSynchronized  ),
            .pe2__sys__ready                            ( pe2__sys__ready             ),
            .pe2__sys__complete                         ( pe2__sys__complete          ),
            // General control and status                  
            .sys__pe3__allSynchronized                  ( sys__pe3__allSynchronized   ),
            .pe3__sys__thisSynchronized                 ( pe3__sys__thisSynchronized  ),
            .pe3__sys__ready                            ( pe3__sys__ready             ),
            .pe3__sys__complete                         ( pe3__sys__complete          ),
            // General control and status                  
            .sys__pe4__allSynchronized                  ( sys__pe4__allSynchronized   ),
            .pe4__sys__thisSynchronized                 ( pe4__sys__thisSynchronized  ),
            .pe4__sys__ready                            ( pe4__sys__ready             ),
            .pe4__sys__complete                         ( pe4__sys__complete          ),
            // General control and status                  
            .sys__pe5__allSynchronized                  ( sys__pe5__allSynchronized   ),
            .pe5__sys__thisSynchronized                 ( pe5__sys__thisSynchronized  ),
            .pe5__sys__ready                            ( pe5__sys__ready             ),
            .pe5__sys__complete                         ( pe5__sys__complete          ),
            // General control and status                  
            .sys__pe6__allSynchronized                  ( sys__pe6__allSynchronized   ),
            .pe6__sys__thisSynchronized                 ( pe6__sys__thisSynchronized  ),
            .pe6__sys__ready                            ( pe6__sys__ready             ),
            .pe6__sys__complete                         ( pe6__sys__complete          ),
            // General control and status                  
            .sys__pe7__allSynchronized                  ( sys__pe7__allSynchronized   ),
            .pe7__sys__thisSynchronized                 ( pe7__sys__thisSynchronized  ),
            .pe7__sys__ready                            ( pe7__sys__ready             ),
            .pe7__sys__complete                         ( pe7__sys__complete          ),
            // General control and status                  
            .sys__pe8__allSynchronized                  ( sys__pe8__allSynchronized   ),
            .pe8__sys__thisSynchronized                 ( pe8__sys__thisSynchronized  ),
            .pe8__sys__ready                            ( pe8__sys__ready             ),
            .pe8__sys__complete                         ( pe8__sys__complete          ),
            // General control and status                  
            .sys__pe9__allSynchronized                  ( sys__pe9__allSynchronized   ),
            .pe9__sys__thisSynchronized                 ( pe9__sys__thisSynchronized  ),
            .pe9__sys__ready                            ( pe9__sys__ready             ),
            .pe9__sys__complete                         ( pe9__sys__complete          ),
            // General control and status                  
            .sys__pe10__allSynchronized                  ( sys__pe10__allSynchronized   ),
            .pe10__sys__thisSynchronized                 ( pe10__sys__thisSynchronized  ),
            .pe10__sys__ready                            ( pe10__sys__ready             ),
            .pe10__sys__complete                         ( pe10__sys__complete          ),
            // General control and status                  
            .sys__pe11__allSynchronized                  ( sys__pe11__allSynchronized   ),
            .pe11__sys__thisSynchronized                 ( pe11__sys__thisSynchronized  ),
            .pe11__sys__ready                            ( pe11__sys__ready             ),
            .pe11__sys__complete                         ( pe11__sys__complete          ),
            // General control and status                  
            .sys__pe12__allSynchronized                  ( sys__pe12__allSynchronized   ),
            .pe12__sys__thisSynchronized                 ( pe12__sys__thisSynchronized  ),
            .pe12__sys__ready                            ( pe12__sys__ready             ),
            .pe12__sys__complete                         ( pe12__sys__complete          ),
            // General control and status                  
            .sys__pe13__allSynchronized                  ( sys__pe13__allSynchronized   ),
            .pe13__sys__thisSynchronized                 ( pe13__sys__thisSynchronized  ),
            .pe13__sys__ready                            ( pe13__sys__ready             ),
            .pe13__sys__complete                         ( pe13__sys__complete          ),
            // General control and status                  
            .sys__pe14__allSynchronized                  ( sys__pe14__allSynchronized   ),
            .pe14__sys__thisSynchronized                 ( pe14__sys__thisSynchronized  ),
            .pe14__sys__ready                            ( pe14__sys__ready             ),
            .pe14__sys__complete                         ( pe14__sys__complete          ),
            // General control and status                  
            .sys__pe15__allSynchronized                  ( sys__pe15__allSynchronized   ),
            .pe15__sys__thisSynchronized                 ( pe15__sys__thisSynchronized  ),
            .pe15__sys__ready                            ( pe15__sys__ready             ),
            .pe15__sys__complete                         ( pe15__sys__complete          ),
            // General control and status                  
            .sys__pe16__allSynchronized                  ( sys__pe16__allSynchronized   ),
            .pe16__sys__thisSynchronized                 ( pe16__sys__thisSynchronized  ),
            .pe16__sys__ready                            ( pe16__sys__ready             ),
            .pe16__sys__complete                         ( pe16__sys__complete          ),
            // General control and status                  
            .sys__pe17__allSynchronized                  ( sys__pe17__allSynchronized   ),
            .pe17__sys__thisSynchronized                 ( pe17__sys__thisSynchronized  ),
            .pe17__sys__ready                            ( pe17__sys__ready             ),
            .pe17__sys__complete                         ( pe17__sys__complete          ),
            // General control and status                  
            .sys__pe18__allSynchronized                  ( sys__pe18__allSynchronized   ),
            .pe18__sys__thisSynchronized                 ( pe18__sys__thisSynchronized  ),
            .pe18__sys__ready                            ( pe18__sys__ready             ),
            .pe18__sys__complete                         ( pe18__sys__complete          ),
            // General control and status                  
            .sys__pe19__allSynchronized                  ( sys__pe19__allSynchronized   ),
            .pe19__sys__thisSynchronized                 ( pe19__sys__thisSynchronized  ),
            .pe19__sys__ready                            ( pe19__sys__ready             ),
            .pe19__sys__complete                         ( pe19__sys__complete          ),
            // General control and status                  
            .sys__pe20__allSynchronized                  ( sys__pe20__allSynchronized   ),
            .pe20__sys__thisSynchronized                 ( pe20__sys__thisSynchronized  ),
            .pe20__sys__ready                            ( pe20__sys__ready             ),
            .pe20__sys__complete                         ( pe20__sys__complete          ),
            // General control and status                  
            .sys__pe21__allSynchronized                  ( sys__pe21__allSynchronized   ),
            .pe21__sys__thisSynchronized                 ( pe21__sys__thisSynchronized  ),
            .pe21__sys__ready                            ( pe21__sys__ready             ),
            .pe21__sys__complete                         ( pe21__sys__complete          ),
            // General control and status                  
            .sys__pe22__allSynchronized                  ( sys__pe22__allSynchronized   ),
            .pe22__sys__thisSynchronized                 ( pe22__sys__thisSynchronized  ),
            .pe22__sys__ready                            ( pe22__sys__ready             ),
            .pe22__sys__complete                         ( pe22__sys__complete          ),
            // General control and status                  
            .sys__pe23__allSynchronized                  ( sys__pe23__allSynchronized   ),
            .pe23__sys__thisSynchronized                 ( pe23__sys__thisSynchronized  ),
            .pe23__sys__ready                            ( pe23__sys__ready             ),
            .pe23__sys__complete                         ( pe23__sys__complete          ),
            // General control and status                  
            .sys__pe24__allSynchronized                  ( sys__pe24__allSynchronized   ),
            .pe24__sys__thisSynchronized                 ( pe24__sys__thisSynchronized  ),
            .pe24__sys__ready                            ( pe24__sys__ready             ),
            .pe24__sys__complete                         ( pe24__sys__complete          ),
            // General control and status                  
            .sys__pe25__allSynchronized                  ( sys__pe25__allSynchronized   ),
            .pe25__sys__thisSynchronized                 ( pe25__sys__thisSynchronized  ),
            .pe25__sys__ready                            ( pe25__sys__ready             ),
            .pe25__sys__complete                         ( pe25__sys__complete          ),
            // General control and status                  
            .sys__pe26__allSynchronized                  ( sys__pe26__allSynchronized   ),
            .pe26__sys__thisSynchronized                 ( pe26__sys__thisSynchronized  ),
            .pe26__sys__ready                            ( pe26__sys__ready             ),
            .pe26__sys__complete                         ( pe26__sys__complete          ),
            // General control and status                  
            .sys__pe27__allSynchronized                  ( sys__pe27__allSynchronized   ),
            .pe27__sys__thisSynchronized                 ( pe27__sys__thisSynchronized  ),
            .pe27__sys__ready                            ( pe27__sys__ready             ),
            .pe27__sys__complete                         ( pe27__sys__complete          ),
            // General control and status                  
            .sys__pe28__allSynchronized                  ( sys__pe28__allSynchronized   ),
            .pe28__sys__thisSynchronized                 ( pe28__sys__thisSynchronized  ),
            .pe28__sys__ready                            ( pe28__sys__ready             ),
            .pe28__sys__complete                         ( pe28__sys__complete          ),
            // General control and status                  
            .sys__pe29__allSynchronized                  ( sys__pe29__allSynchronized   ),
            .pe29__sys__thisSynchronized                 ( pe29__sys__thisSynchronized  ),
            .pe29__sys__ready                            ( pe29__sys__ready             ),
            .pe29__sys__complete                         ( pe29__sys__complete          ),
            // General control and status                  
            .sys__pe30__allSynchronized                  ( sys__pe30__allSynchronized   ),
            .pe30__sys__thisSynchronized                 ( pe30__sys__thisSynchronized  ),
            .pe30__sys__ready                            ( pe30__sys__ready             ),
            .pe30__sys__complete                         ( pe30__sys__complete          ),
            // General control and status                  
            .sys__pe31__allSynchronized                  ( sys__pe31__allSynchronized   ),
            .pe31__sys__thisSynchronized                 ( pe31__sys__thisSynchronized  ),
            .pe31__sys__ready                            ( pe31__sys__ready             ),
            .pe31__sys__complete                         ( pe31__sys__complete          ),
            // General control and status                  
            .sys__pe32__allSynchronized                  ( sys__pe32__allSynchronized   ),
            .pe32__sys__thisSynchronized                 ( pe32__sys__thisSynchronized  ),
            .pe32__sys__ready                            ( pe32__sys__ready             ),
            .pe32__sys__complete                         ( pe32__sys__complete          ),
            // General control and status                  
            .sys__pe33__allSynchronized                  ( sys__pe33__allSynchronized   ),
            .pe33__sys__thisSynchronized                 ( pe33__sys__thisSynchronized  ),
            .pe33__sys__ready                            ( pe33__sys__ready             ),
            .pe33__sys__complete                         ( pe33__sys__complete          ),
            // General control and status                  
            .sys__pe34__allSynchronized                  ( sys__pe34__allSynchronized   ),
            .pe34__sys__thisSynchronized                 ( pe34__sys__thisSynchronized  ),
            .pe34__sys__ready                            ( pe34__sys__ready             ),
            .pe34__sys__complete                         ( pe34__sys__complete          ),
            // General control and status                  
            .sys__pe35__allSynchronized                  ( sys__pe35__allSynchronized   ),
            .pe35__sys__thisSynchronized                 ( pe35__sys__thisSynchronized  ),
            .pe35__sys__ready                            ( pe35__sys__ready             ),
            .pe35__sys__complete                         ( pe35__sys__complete          ),
            // General control and status                  
            .sys__pe36__allSynchronized                  ( sys__pe36__allSynchronized   ),
            .pe36__sys__thisSynchronized                 ( pe36__sys__thisSynchronized  ),
            .pe36__sys__ready                            ( pe36__sys__ready             ),
            .pe36__sys__complete                         ( pe36__sys__complete          ),
            // General control and status                  
            .sys__pe37__allSynchronized                  ( sys__pe37__allSynchronized   ),
            .pe37__sys__thisSynchronized                 ( pe37__sys__thisSynchronized  ),
            .pe37__sys__ready                            ( pe37__sys__ready             ),
            .pe37__sys__complete                         ( pe37__sys__complete          ),
            // General control and status                  
            .sys__pe38__allSynchronized                  ( sys__pe38__allSynchronized   ),
            .pe38__sys__thisSynchronized                 ( pe38__sys__thisSynchronized  ),
            .pe38__sys__ready                            ( pe38__sys__ready             ),
            .pe38__sys__complete                         ( pe38__sys__complete          ),
            // General control and status                  
            .sys__pe39__allSynchronized                  ( sys__pe39__allSynchronized   ),
            .pe39__sys__thisSynchronized                 ( pe39__sys__thisSynchronized  ),
            .pe39__sys__ready                            ( pe39__sys__ready             ),
            .pe39__sys__complete                         ( pe39__sys__complete          ),
            // General control and status                  
            .sys__pe40__allSynchronized                  ( sys__pe40__allSynchronized   ),
            .pe40__sys__thisSynchronized                 ( pe40__sys__thisSynchronized  ),
            .pe40__sys__ready                            ( pe40__sys__ready             ),
            .pe40__sys__complete                         ( pe40__sys__complete          ),
            // General control and status                  
            .sys__pe41__allSynchronized                  ( sys__pe41__allSynchronized   ),
            .pe41__sys__thisSynchronized                 ( pe41__sys__thisSynchronized  ),
            .pe41__sys__ready                            ( pe41__sys__ready             ),
            .pe41__sys__complete                         ( pe41__sys__complete          ),
            // General control and status                  
            .sys__pe42__allSynchronized                  ( sys__pe42__allSynchronized   ),
            .pe42__sys__thisSynchronized                 ( pe42__sys__thisSynchronized  ),
            .pe42__sys__ready                            ( pe42__sys__ready             ),
            .pe42__sys__complete                         ( pe42__sys__complete          ),
            // General control and status                  
            .sys__pe43__allSynchronized                  ( sys__pe43__allSynchronized   ),
            .pe43__sys__thisSynchronized                 ( pe43__sys__thisSynchronized  ),
            .pe43__sys__ready                            ( pe43__sys__ready             ),
            .pe43__sys__complete                         ( pe43__sys__complete          ),
            // General control and status                  
            .sys__pe44__allSynchronized                  ( sys__pe44__allSynchronized   ),
            .pe44__sys__thisSynchronized                 ( pe44__sys__thisSynchronized  ),
            .pe44__sys__ready                            ( pe44__sys__ready             ),
            .pe44__sys__complete                         ( pe44__sys__complete          ),
            // General control and status                  
            .sys__pe45__allSynchronized                  ( sys__pe45__allSynchronized   ),
            .pe45__sys__thisSynchronized                 ( pe45__sys__thisSynchronized  ),
            .pe45__sys__ready                            ( pe45__sys__ready             ),
            .pe45__sys__complete                         ( pe45__sys__complete          ),
            // General control and status                  
            .sys__pe46__allSynchronized                  ( sys__pe46__allSynchronized   ),
            .pe46__sys__thisSynchronized                 ( pe46__sys__thisSynchronized  ),
            .pe46__sys__ready                            ( pe46__sys__ready             ),
            .pe46__sys__complete                         ( pe46__sys__complete          ),
            // General control and status                  
            .sys__pe47__allSynchronized                  ( sys__pe47__allSynchronized   ),
            .pe47__sys__thisSynchronized                 ( pe47__sys__thisSynchronized  ),
            .pe47__sys__ready                            ( pe47__sys__ready             ),
            .pe47__sys__complete                         ( pe47__sys__complete          ),
            // General control and status                  
            .sys__pe48__allSynchronized                  ( sys__pe48__allSynchronized   ),
            .pe48__sys__thisSynchronized                 ( pe48__sys__thisSynchronized  ),
            .pe48__sys__ready                            ( pe48__sys__ready             ),
            .pe48__sys__complete                         ( pe48__sys__complete          ),
            // General control and status                  
            .sys__pe49__allSynchronized                  ( sys__pe49__allSynchronized   ),
            .pe49__sys__thisSynchronized                 ( pe49__sys__thisSynchronized  ),
            .pe49__sys__ready                            ( pe49__sys__ready             ),
            .pe49__sys__complete                         ( pe49__sys__complete          ),
            // General control and status                  
            .sys__pe50__allSynchronized                  ( sys__pe50__allSynchronized   ),
            .pe50__sys__thisSynchronized                 ( pe50__sys__thisSynchronized  ),
            .pe50__sys__ready                            ( pe50__sys__ready             ),
            .pe50__sys__complete                         ( pe50__sys__complete          ),
            // General control and status                  
            .sys__pe51__allSynchronized                  ( sys__pe51__allSynchronized   ),
            .pe51__sys__thisSynchronized                 ( pe51__sys__thisSynchronized  ),
            .pe51__sys__ready                            ( pe51__sys__ready             ),
            .pe51__sys__complete                         ( pe51__sys__complete          ),
            // General control and status                  
            .sys__pe52__allSynchronized                  ( sys__pe52__allSynchronized   ),
            .pe52__sys__thisSynchronized                 ( pe52__sys__thisSynchronized  ),
            .pe52__sys__ready                            ( pe52__sys__ready             ),
            .pe52__sys__complete                         ( pe52__sys__complete          ),
            // General control and status                  
            .sys__pe53__allSynchronized                  ( sys__pe53__allSynchronized   ),
            .pe53__sys__thisSynchronized                 ( pe53__sys__thisSynchronized  ),
            .pe53__sys__ready                            ( pe53__sys__ready             ),
            .pe53__sys__complete                         ( pe53__sys__complete          ),
            // General control and status                  
            .sys__pe54__allSynchronized                  ( sys__pe54__allSynchronized   ),
            .pe54__sys__thisSynchronized                 ( pe54__sys__thisSynchronized  ),
            .pe54__sys__ready                            ( pe54__sys__ready             ),
            .pe54__sys__complete                         ( pe54__sys__complete          ),
            // General control and status                  
            .sys__pe55__allSynchronized                  ( sys__pe55__allSynchronized   ),
            .pe55__sys__thisSynchronized                 ( pe55__sys__thisSynchronized  ),
            .pe55__sys__ready                            ( pe55__sys__ready             ),
            .pe55__sys__complete                         ( pe55__sys__complete          ),
            // General control and status                  
            .sys__pe56__allSynchronized                  ( sys__pe56__allSynchronized   ),
            .pe56__sys__thisSynchronized                 ( pe56__sys__thisSynchronized  ),
            .pe56__sys__ready                            ( pe56__sys__ready             ),
            .pe56__sys__complete                         ( pe56__sys__complete          ),
            // General control and status                  
            .sys__pe57__allSynchronized                  ( sys__pe57__allSynchronized   ),
            .pe57__sys__thisSynchronized                 ( pe57__sys__thisSynchronized  ),
            .pe57__sys__ready                            ( pe57__sys__ready             ),
            .pe57__sys__complete                         ( pe57__sys__complete          ),
            // General control and status                  
            .sys__pe58__allSynchronized                  ( sys__pe58__allSynchronized   ),
            .pe58__sys__thisSynchronized                 ( pe58__sys__thisSynchronized  ),
            .pe58__sys__ready                            ( pe58__sys__ready             ),
            .pe58__sys__complete                         ( pe58__sys__complete          ),
            // General control and status                  
            .sys__pe59__allSynchronized                  ( sys__pe59__allSynchronized   ),
            .pe59__sys__thisSynchronized                 ( pe59__sys__thisSynchronized  ),
            .pe59__sys__ready                            ( pe59__sys__ready             ),
            .pe59__sys__complete                         ( pe59__sys__complete          ),
            // General control and status                  
            .sys__pe60__allSynchronized                  ( sys__pe60__allSynchronized   ),
            .pe60__sys__thisSynchronized                 ( pe60__sys__thisSynchronized  ),
            .pe60__sys__ready                            ( pe60__sys__ready             ),
            .pe60__sys__complete                         ( pe60__sys__complete          ),
            // General control and status                  
            .sys__pe61__allSynchronized                  ( sys__pe61__allSynchronized   ),
            .pe61__sys__thisSynchronized                 ( pe61__sys__thisSynchronized  ),
            .pe61__sys__ready                            ( pe61__sys__ready             ),
            .pe61__sys__complete                         ( pe61__sys__complete          ),
            // General control and status                  
            .sys__pe62__allSynchronized                  ( sys__pe62__allSynchronized   ),
            .pe62__sys__thisSynchronized                 ( pe62__sys__thisSynchronized  ),
            .pe62__sys__ready                            ( pe62__sys__ready             ),
            .pe62__sys__complete                         ( pe62__sys__complete          ),
            // General control and status                  
            .sys__pe63__allSynchronized                  ( sys__pe63__allSynchronized   ),
            .pe63__sys__thisSynchronized                 ( pe63__sys__thisSynchronized  ),
            .pe63__sys__ready                            ( pe63__sys__ready             ),
            .pe63__sys__complete                         ( pe63__sys__complete          ),