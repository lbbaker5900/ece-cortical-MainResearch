
  reg [31:0] pe0_lane0_strm0 [0:4095];
  reg [31:0] pe0_lane0_strm0_tmp     ;
  reg [31:0] pe0_lane0_strm1 [0:4095];
  reg [31:0] pe0_lane0_strm1_tmp     ;
  reg [31:0] pe0_lane1_strm0 [0:4095];
  reg [31:0] pe0_lane1_strm0_tmp     ;
  reg [31:0] pe0_lane1_strm1 [0:4095];
  reg [31:0] pe0_lane1_strm1_tmp     ;
  reg [31:0] pe0_lane2_strm0 [0:4095];
  reg [31:0] pe0_lane2_strm0_tmp     ;
  reg [31:0] pe0_lane2_strm1 [0:4095];
  reg [31:0] pe0_lane2_strm1_tmp     ;
  reg [31:0] pe0_lane3_strm0 [0:4095];
  reg [31:0] pe0_lane3_strm0_tmp     ;
  reg [31:0] pe0_lane3_strm1 [0:4095];
  reg [31:0] pe0_lane3_strm1_tmp     ;
  reg [31:0] pe0_lane4_strm0 [0:4095];
  reg [31:0] pe0_lane4_strm0_tmp     ;
  reg [31:0] pe0_lane4_strm1 [0:4095];
  reg [31:0] pe0_lane4_strm1_tmp     ;
  reg [31:0] pe0_lane5_strm0 [0:4095];
  reg [31:0] pe0_lane5_strm0_tmp     ;
  reg [31:0] pe0_lane5_strm1 [0:4095];
  reg [31:0] pe0_lane5_strm1_tmp     ;
  reg [31:0] pe0_lane6_strm0 [0:4095];
  reg [31:0] pe0_lane6_strm0_tmp     ;
  reg [31:0] pe0_lane6_strm1 [0:4095];
  reg [31:0] pe0_lane6_strm1_tmp     ;
  reg [31:0] pe0_lane7_strm0 [0:4095];
  reg [31:0] pe0_lane7_strm0_tmp     ;
  reg [31:0] pe0_lane7_strm1 [0:4095];
  reg [31:0] pe0_lane7_strm1_tmp     ;
  reg [31:0] pe0_lane8_strm0 [0:4095];
  reg [31:0] pe0_lane8_strm0_tmp     ;
  reg [31:0] pe0_lane8_strm1 [0:4095];
  reg [31:0] pe0_lane8_strm1_tmp     ;
  reg [31:0] pe0_lane9_strm0 [0:4095];
  reg [31:0] pe0_lane9_strm0_tmp     ;
  reg [31:0] pe0_lane9_strm1 [0:4095];
  reg [31:0] pe0_lane9_strm1_tmp     ;
  reg [31:0] pe0_lane10_strm0 [0:4095];
  reg [31:0] pe0_lane10_strm0_tmp     ;
  reg [31:0] pe0_lane10_strm1 [0:4095];
  reg [31:0] pe0_lane10_strm1_tmp     ;
  reg [31:0] pe0_lane11_strm0 [0:4095];
  reg [31:0] pe0_lane11_strm0_tmp     ;
  reg [31:0] pe0_lane11_strm1 [0:4095];
  reg [31:0] pe0_lane11_strm1_tmp     ;
  reg [31:0] pe0_lane12_strm0 [0:4095];
  reg [31:0] pe0_lane12_strm0_tmp     ;
  reg [31:0] pe0_lane12_strm1 [0:4095];
  reg [31:0] pe0_lane12_strm1_tmp     ;
  reg [31:0] pe0_lane13_strm0 [0:4095];
  reg [31:0] pe0_lane13_strm0_tmp     ;
  reg [31:0] pe0_lane13_strm1 [0:4095];
  reg [31:0] pe0_lane13_strm1_tmp     ;
  reg [31:0] pe0_lane14_strm0 [0:4095];
  reg [31:0] pe0_lane14_strm0_tmp     ;
  reg [31:0] pe0_lane14_strm1 [0:4095];
  reg [31:0] pe0_lane14_strm1_tmp     ;
  reg [31:0] pe0_lane15_strm0 [0:4095];
  reg [31:0] pe0_lane15_strm0_tmp     ;
  reg [31:0] pe0_lane15_strm1 [0:4095];
  reg [31:0] pe0_lane15_strm1_tmp     ;
  reg [31:0] pe0_lane16_strm0 [0:4095];
  reg [31:0] pe0_lane16_strm0_tmp     ;
  reg [31:0] pe0_lane16_strm1 [0:4095];
  reg [31:0] pe0_lane16_strm1_tmp     ;
  reg [31:0] pe0_lane17_strm0 [0:4095];
  reg [31:0] pe0_lane17_strm0_tmp     ;
  reg [31:0] pe0_lane17_strm1 [0:4095];
  reg [31:0] pe0_lane17_strm1_tmp     ;
  reg [31:0] pe0_lane18_strm0 [0:4095];
  reg [31:0] pe0_lane18_strm0_tmp     ;
  reg [31:0] pe0_lane18_strm1 [0:4095];
  reg [31:0] pe0_lane18_strm1_tmp     ;
  reg [31:0] pe0_lane19_strm0 [0:4095];
  reg [31:0] pe0_lane19_strm0_tmp     ;
  reg [31:0] pe0_lane19_strm1 [0:4095];
  reg [31:0] pe0_lane19_strm1_tmp     ;
  reg [31:0] pe0_lane20_strm0 [0:4095];
  reg [31:0] pe0_lane20_strm0_tmp     ;
  reg [31:0] pe0_lane20_strm1 [0:4095];
  reg [31:0] pe0_lane20_strm1_tmp     ;
  reg [31:0] pe0_lane21_strm0 [0:4095];
  reg [31:0] pe0_lane21_strm0_tmp     ;
  reg [31:0] pe0_lane21_strm1 [0:4095];
  reg [31:0] pe0_lane21_strm1_tmp     ;
  reg [31:0] pe0_lane22_strm0 [0:4095];
  reg [31:0] pe0_lane22_strm0_tmp     ;
  reg [31:0] pe0_lane22_strm1 [0:4095];
  reg [31:0] pe0_lane22_strm1_tmp     ;
  reg [31:0] pe0_lane23_strm0 [0:4095];
  reg [31:0] pe0_lane23_strm0_tmp     ;
  reg [31:0] pe0_lane23_strm1 [0:4095];
  reg [31:0] pe0_lane23_strm1_tmp     ;
  reg [31:0] pe0_lane24_strm0 [0:4095];
  reg [31:0] pe0_lane24_strm0_tmp     ;
  reg [31:0] pe0_lane24_strm1 [0:4095];
  reg [31:0] pe0_lane24_strm1_tmp     ;
  reg [31:0] pe0_lane25_strm0 [0:4095];
  reg [31:0] pe0_lane25_strm0_tmp     ;
  reg [31:0] pe0_lane25_strm1 [0:4095];
  reg [31:0] pe0_lane25_strm1_tmp     ;
  reg [31:0] pe0_lane26_strm0 [0:4095];
  reg [31:0] pe0_lane26_strm0_tmp     ;
  reg [31:0] pe0_lane26_strm1 [0:4095];
  reg [31:0] pe0_lane26_strm1_tmp     ;
  reg [31:0] pe0_lane27_strm0 [0:4095];
  reg [31:0] pe0_lane27_strm0_tmp     ;
  reg [31:0] pe0_lane27_strm1 [0:4095];
  reg [31:0] pe0_lane27_strm1_tmp     ;
  reg [31:0] pe0_lane28_strm0 [0:4095];
  reg [31:0] pe0_lane28_strm0_tmp     ;
  reg [31:0] pe0_lane28_strm1 [0:4095];
  reg [31:0] pe0_lane28_strm1_tmp     ;
  reg [31:0] pe0_lane29_strm0 [0:4095];
  reg [31:0] pe0_lane29_strm0_tmp     ;
  reg [31:0] pe0_lane29_strm1 [0:4095];
  reg [31:0] pe0_lane29_strm1_tmp     ;
  reg [31:0] pe0_lane30_strm0 [0:4095];
  reg [31:0] pe0_lane30_strm0_tmp     ;
  reg [31:0] pe0_lane30_strm1 [0:4095];
  reg [31:0] pe0_lane30_strm1_tmp     ;
  reg [31:0] pe0_lane31_strm0 [0:4095];
  reg [31:0] pe0_lane31_strm0_tmp     ;
  reg [31:0] pe0_lane31_strm1 [0:4095];
  reg [31:0] pe0_lane31_strm1_tmp     ;
  reg [31:0] pe1_lane0_strm0 [0:4095];
  reg [31:0] pe1_lane0_strm0_tmp     ;
  reg [31:0] pe1_lane0_strm1 [0:4095];
  reg [31:0] pe1_lane0_strm1_tmp     ;
  reg [31:0] pe1_lane1_strm0 [0:4095];
  reg [31:0] pe1_lane1_strm0_tmp     ;
  reg [31:0] pe1_lane1_strm1 [0:4095];
  reg [31:0] pe1_lane1_strm1_tmp     ;
  reg [31:0] pe1_lane2_strm0 [0:4095];
  reg [31:0] pe1_lane2_strm0_tmp     ;
  reg [31:0] pe1_lane2_strm1 [0:4095];
  reg [31:0] pe1_lane2_strm1_tmp     ;
  reg [31:0] pe1_lane3_strm0 [0:4095];
  reg [31:0] pe1_lane3_strm0_tmp     ;
  reg [31:0] pe1_lane3_strm1 [0:4095];
  reg [31:0] pe1_lane3_strm1_tmp     ;
  reg [31:0] pe1_lane4_strm0 [0:4095];
  reg [31:0] pe1_lane4_strm0_tmp     ;
  reg [31:0] pe1_lane4_strm1 [0:4095];
  reg [31:0] pe1_lane4_strm1_tmp     ;
  reg [31:0] pe1_lane5_strm0 [0:4095];
  reg [31:0] pe1_lane5_strm0_tmp     ;
  reg [31:0] pe1_lane5_strm1 [0:4095];
  reg [31:0] pe1_lane5_strm1_tmp     ;
  reg [31:0] pe1_lane6_strm0 [0:4095];
  reg [31:0] pe1_lane6_strm0_tmp     ;
  reg [31:0] pe1_lane6_strm1 [0:4095];
  reg [31:0] pe1_lane6_strm1_tmp     ;
  reg [31:0] pe1_lane7_strm0 [0:4095];
  reg [31:0] pe1_lane7_strm0_tmp     ;
  reg [31:0] pe1_lane7_strm1 [0:4095];
  reg [31:0] pe1_lane7_strm1_tmp     ;
  reg [31:0] pe1_lane8_strm0 [0:4095];
  reg [31:0] pe1_lane8_strm0_tmp     ;
  reg [31:0] pe1_lane8_strm1 [0:4095];
  reg [31:0] pe1_lane8_strm1_tmp     ;
  reg [31:0] pe1_lane9_strm0 [0:4095];
  reg [31:0] pe1_lane9_strm0_tmp     ;
  reg [31:0] pe1_lane9_strm1 [0:4095];
  reg [31:0] pe1_lane9_strm1_tmp     ;
  reg [31:0] pe1_lane10_strm0 [0:4095];
  reg [31:0] pe1_lane10_strm0_tmp     ;
  reg [31:0] pe1_lane10_strm1 [0:4095];
  reg [31:0] pe1_lane10_strm1_tmp     ;
  reg [31:0] pe1_lane11_strm0 [0:4095];
  reg [31:0] pe1_lane11_strm0_tmp     ;
  reg [31:0] pe1_lane11_strm1 [0:4095];
  reg [31:0] pe1_lane11_strm1_tmp     ;
  reg [31:0] pe1_lane12_strm0 [0:4095];
  reg [31:0] pe1_lane12_strm0_tmp     ;
  reg [31:0] pe1_lane12_strm1 [0:4095];
  reg [31:0] pe1_lane12_strm1_tmp     ;
  reg [31:0] pe1_lane13_strm0 [0:4095];
  reg [31:0] pe1_lane13_strm0_tmp     ;
  reg [31:0] pe1_lane13_strm1 [0:4095];
  reg [31:0] pe1_lane13_strm1_tmp     ;
  reg [31:0] pe1_lane14_strm0 [0:4095];
  reg [31:0] pe1_lane14_strm0_tmp     ;
  reg [31:0] pe1_lane14_strm1 [0:4095];
  reg [31:0] pe1_lane14_strm1_tmp     ;
  reg [31:0] pe1_lane15_strm0 [0:4095];
  reg [31:0] pe1_lane15_strm0_tmp     ;
  reg [31:0] pe1_lane15_strm1 [0:4095];
  reg [31:0] pe1_lane15_strm1_tmp     ;
  reg [31:0] pe1_lane16_strm0 [0:4095];
  reg [31:0] pe1_lane16_strm0_tmp     ;
  reg [31:0] pe1_lane16_strm1 [0:4095];
  reg [31:0] pe1_lane16_strm1_tmp     ;
  reg [31:0] pe1_lane17_strm0 [0:4095];
  reg [31:0] pe1_lane17_strm0_tmp     ;
  reg [31:0] pe1_lane17_strm1 [0:4095];
  reg [31:0] pe1_lane17_strm1_tmp     ;
  reg [31:0] pe1_lane18_strm0 [0:4095];
  reg [31:0] pe1_lane18_strm0_tmp     ;
  reg [31:0] pe1_lane18_strm1 [0:4095];
  reg [31:0] pe1_lane18_strm1_tmp     ;
  reg [31:0] pe1_lane19_strm0 [0:4095];
  reg [31:0] pe1_lane19_strm0_tmp     ;
  reg [31:0] pe1_lane19_strm1 [0:4095];
  reg [31:0] pe1_lane19_strm1_tmp     ;
  reg [31:0] pe1_lane20_strm0 [0:4095];
  reg [31:0] pe1_lane20_strm0_tmp     ;
  reg [31:0] pe1_lane20_strm1 [0:4095];
  reg [31:0] pe1_lane20_strm1_tmp     ;
  reg [31:0] pe1_lane21_strm0 [0:4095];
  reg [31:0] pe1_lane21_strm0_tmp     ;
  reg [31:0] pe1_lane21_strm1 [0:4095];
  reg [31:0] pe1_lane21_strm1_tmp     ;
  reg [31:0] pe1_lane22_strm0 [0:4095];
  reg [31:0] pe1_lane22_strm0_tmp     ;
  reg [31:0] pe1_lane22_strm1 [0:4095];
  reg [31:0] pe1_lane22_strm1_tmp     ;
  reg [31:0] pe1_lane23_strm0 [0:4095];
  reg [31:0] pe1_lane23_strm0_tmp     ;
  reg [31:0] pe1_lane23_strm1 [0:4095];
  reg [31:0] pe1_lane23_strm1_tmp     ;
  reg [31:0] pe1_lane24_strm0 [0:4095];
  reg [31:0] pe1_lane24_strm0_tmp     ;
  reg [31:0] pe1_lane24_strm1 [0:4095];
  reg [31:0] pe1_lane24_strm1_tmp     ;
  reg [31:0] pe1_lane25_strm0 [0:4095];
  reg [31:0] pe1_lane25_strm0_tmp     ;
  reg [31:0] pe1_lane25_strm1 [0:4095];
  reg [31:0] pe1_lane25_strm1_tmp     ;
  reg [31:0] pe1_lane26_strm0 [0:4095];
  reg [31:0] pe1_lane26_strm0_tmp     ;
  reg [31:0] pe1_lane26_strm1 [0:4095];
  reg [31:0] pe1_lane26_strm1_tmp     ;
  reg [31:0] pe1_lane27_strm0 [0:4095];
  reg [31:0] pe1_lane27_strm0_tmp     ;
  reg [31:0] pe1_lane27_strm1 [0:4095];
  reg [31:0] pe1_lane27_strm1_tmp     ;
  reg [31:0] pe1_lane28_strm0 [0:4095];
  reg [31:0] pe1_lane28_strm0_tmp     ;
  reg [31:0] pe1_lane28_strm1 [0:4095];
  reg [31:0] pe1_lane28_strm1_tmp     ;
  reg [31:0] pe1_lane29_strm0 [0:4095];
  reg [31:0] pe1_lane29_strm0_tmp     ;
  reg [31:0] pe1_lane29_strm1 [0:4095];
  reg [31:0] pe1_lane29_strm1_tmp     ;
  reg [31:0] pe1_lane30_strm0 [0:4095];
  reg [31:0] pe1_lane30_strm0_tmp     ;
  reg [31:0] pe1_lane30_strm1 [0:4095];
  reg [31:0] pe1_lane30_strm1_tmp     ;
  reg [31:0] pe1_lane31_strm0 [0:4095];
  reg [31:0] pe1_lane31_strm0_tmp     ;
  reg [31:0] pe1_lane31_strm1 [0:4095];
  reg [31:0] pe1_lane31_strm1_tmp     ;
  reg [31:0] pe2_lane0_strm0 [0:4095];
  reg [31:0] pe2_lane0_strm0_tmp     ;
  reg [31:0] pe2_lane0_strm1 [0:4095];
  reg [31:0] pe2_lane0_strm1_tmp     ;
  reg [31:0] pe2_lane1_strm0 [0:4095];
  reg [31:0] pe2_lane1_strm0_tmp     ;
  reg [31:0] pe2_lane1_strm1 [0:4095];
  reg [31:0] pe2_lane1_strm1_tmp     ;
  reg [31:0] pe2_lane2_strm0 [0:4095];
  reg [31:0] pe2_lane2_strm0_tmp     ;
  reg [31:0] pe2_lane2_strm1 [0:4095];
  reg [31:0] pe2_lane2_strm1_tmp     ;
  reg [31:0] pe2_lane3_strm0 [0:4095];
  reg [31:0] pe2_lane3_strm0_tmp     ;
  reg [31:0] pe2_lane3_strm1 [0:4095];
  reg [31:0] pe2_lane3_strm1_tmp     ;
  reg [31:0] pe2_lane4_strm0 [0:4095];
  reg [31:0] pe2_lane4_strm0_tmp     ;
  reg [31:0] pe2_lane4_strm1 [0:4095];
  reg [31:0] pe2_lane4_strm1_tmp     ;
  reg [31:0] pe2_lane5_strm0 [0:4095];
  reg [31:0] pe2_lane5_strm0_tmp     ;
  reg [31:0] pe2_lane5_strm1 [0:4095];
  reg [31:0] pe2_lane5_strm1_tmp     ;
  reg [31:0] pe2_lane6_strm0 [0:4095];
  reg [31:0] pe2_lane6_strm0_tmp     ;
  reg [31:0] pe2_lane6_strm1 [0:4095];
  reg [31:0] pe2_lane6_strm1_tmp     ;
  reg [31:0] pe2_lane7_strm0 [0:4095];
  reg [31:0] pe2_lane7_strm0_tmp     ;
  reg [31:0] pe2_lane7_strm1 [0:4095];
  reg [31:0] pe2_lane7_strm1_tmp     ;
  reg [31:0] pe2_lane8_strm0 [0:4095];
  reg [31:0] pe2_lane8_strm0_tmp     ;
  reg [31:0] pe2_lane8_strm1 [0:4095];
  reg [31:0] pe2_lane8_strm1_tmp     ;
  reg [31:0] pe2_lane9_strm0 [0:4095];
  reg [31:0] pe2_lane9_strm0_tmp     ;
  reg [31:0] pe2_lane9_strm1 [0:4095];
  reg [31:0] pe2_lane9_strm1_tmp     ;
  reg [31:0] pe2_lane10_strm0 [0:4095];
  reg [31:0] pe2_lane10_strm0_tmp     ;
  reg [31:0] pe2_lane10_strm1 [0:4095];
  reg [31:0] pe2_lane10_strm1_tmp     ;
  reg [31:0] pe2_lane11_strm0 [0:4095];
  reg [31:0] pe2_lane11_strm0_tmp     ;
  reg [31:0] pe2_lane11_strm1 [0:4095];
  reg [31:0] pe2_lane11_strm1_tmp     ;
  reg [31:0] pe2_lane12_strm0 [0:4095];
  reg [31:0] pe2_lane12_strm0_tmp     ;
  reg [31:0] pe2_lane12_strm1 [0:4095];
  reg [31:0] pe2_lane12_strm1_tmp     ;
  reg [31:0] pe2_lane13_strm0 [0:4095];
  reg [31:0] pe2_lane13_strm0_tmp     ;
  reg [31:0] pe2_lane13_strm1 [0:4095];
  reg [31:0] pe2_lane13_strm1_tmp     ;
  reg [31:0] pe2_lane14_strm0 [0:4095];
  reg [31:0] pe2_lane14_strm0_tmp     ;
  reg [31:0] pe2_lane14_strm1 [0:4095];
  reg [31:0] pe2_lane14_strm1_tmp     ;
  reg [31:0] pe2_lane15_strm0 [0:4095];
  reg [31:0] pe2_lane15_strm0_tmp     ;
  reg [31:0] pe2_lane15_strm1 [0:4095];
  reg [31:0] pe2_lane15_strm1_tmp     ;
  reg [31:0] pe2_lane16_strm0 [0:4095];
  reg [31:0] pe2_lane16_strm0_tmp     ;
  reg [31:0] pe2_lane16_strm1 [0:4095];
  reg [31:0] pe2_lane16_strm1_tmp     ;
  reg [31:0] pe2_lane17_strm0 [0:4095];
  reg [31:0] pe2_lane17_strm0_tmp     ;
  reg [31:0] pe2_lane17_strm1 [0:4095];
  reg [31:0] pe2_lane17_strm1_tmp     ;
  reg [31:0] pe2_lane18_strm0 [0:4095];
  reg [31:0] pe2_lane18_strm0_tmp     ;
  reg [31:0] pe2_lane18_strm1 [0:4095];
  reg [31:0] pe2_lane18_strm1_tmp     ;
  reg [31:0] pe2_lane19_strm0 [0:4095];
  reg [31:0] pe2_lane19_strm0_tmp     ;
  reg [31:0] pe2_lane19_strm1 [0:4095];
  reg [31:0] pe2_lane19_strm1_tmp     ;
  reg [31:0] pe2_lane20_strm0 [0:4095];
  reg [31:0] pe2_lane20_strm0_tmp     ;
  reg [31:0] pe2_lane20_strm1 [0:4095];
  reg [31:0] pe2_lane20_strm1_tmp     ;
  reg [31:0] pe2_lane21_strm0 [0:4095];
  reg [31:0] pe2_lane21_strm0_tmp     ;
  reg [31:0] pe2_lane21_strm1 [0:4095];
  reg [31:0] pe2_lane21_strm1_tmp     ;
  reg [31:0] pe2_lane22_strm0 [0:4095];
  reg [31:0] pe2_lane22_strm0_tmp     ;
  reg [31:0] pe2_lane22_strm1 [0:4095];
  reg [31:0] pe2_lane22_strm1_tmp     ;
  reg [31:0] pe2_lane23_strm0 [0:4095];
  reg [31:0] pe2_lane23_strm0_tmp     ;
  reg [31:0] pe2_lane23_strm1 [0:4095];
  reg [31:0] pe2_lane23_strm1_tmp     ;
  reg [31:0] pe2_lane24_strm0 [0:4095];
  reg [31:0] pe2_lane24_strm0_tmp     ;
  reg [31:0] pe2_lane24_strm1 [0:4095];
  reg [31:0] pe2_lane24_strm1_tmp     ;
  reg [31:0] pe2_lane25_strm0 [0:4095];
  reg [31:0] pe2_lane25_strm0_tmp     ;
  reg [31:0] pe2_lane25_strm1 [0:4095];
  reg [31:0] pe2_lane25_strm1_tmp     ;
  reg [31:0] pe2_lane26_strm0 [0:4095];
  reg [31:0] pe2_lane26_strm0_tmp     ;
  reg [31:0] pe2_lane26_strm1 [0:4095];
  reg [31:0] pe2_lane26_strm1_tmp     ;
  reg [31:0] pe2_lane27_strm0 [0:4095];
  reg [31:0] pe2_lane27_strm0_tmp     ;
  reg [31:0] pe2_lane27_strm1 [0:4095];
  reg [31:0] pe2_lane27_strm1_tmp     ;
  reg [31:0] pe2_lane28_strm0 [0:4095];
  reg [31:0] pe2_lane28_strm0_tmp     ;
  reg [31:0] pe2_lane28_strm1 [0:4095];
  reg [31:0] pe2_lane28_strm1_tmp     ;
  reg [31:0] pe2_lane29_strm0 [0:4095];
  reg [31:0] pe2_lane29_strm0_tmp     ;
  reg [31:0] pe2_lane29_strm1 [0:4095];
  reg [31:0] pe2_lane29_strm1_tmp     ;
  reg [31:0] pe2_lane30_strm0 [0:4095];
  reg [31:0] pe2_lane30_strm0_tmp     ;
  reg [31:0] pe2_lane30_strm1 [0:4095];
  reg [31:0] pe2_lane30_strm1_tmp     ;
  reg [31:0] pe2_lane31_strm0 [0:4095];
  reg [31:0] pe2_lane31_strm0_tmp     ;
  reg [31:0] pe2_lane31_strm1 [0:4095];
  reg [31:0] pe2_lane31_strm1_tmp     ;
  reg [31:0] pe3_lane0_strm0 [0:4095];
  reg [31:0] pe3_lane0_strm0_tmp     ;
  reg [31:0] pe3_lane0_strm1 [0:4095];
  reg [31:0] pe3_lane0_strm1_tmp     ;
  reg [31:0] pe3_lane1_strm0 [0:4095];
  reg [31:0] pe3_lane1_strm0_tmp     ;
  reg [31:0] pe3_lane1_strm1 [0:4095];
  reg [31:0] pe3_lane1_strm1_tmp     ;
  reg [31:0] pe3_lane2_strm0 [0:4095];
  reg [31:0] pe3_lane2_strm0_tmp     ;
  reg [31:0] pe3_lane2_strm1 [0:4095];
  reg [31:0] pe3_lane2_strm1_tmp     ;
  reg [31:0] pe3_lane3_strm0 [0:4095];
  reg [31:0] pe3_lane3_strm0_tmp     ;
  reg [31:0] pe3_lane3_strm1 [0:4095];
  reg [31:0] pe3_lane3_strm1_tmp     ;
  reg [31:0] pe3_lane4_strm0 [0:4095];
  reg [31:0] pe3_lane4_strm0_tmp     ;
  reg [31:0] pe3_lane4_strm1 [0:4095];
  reg [31:0] pe3_lane4_strm1_tmp     ;
  reg [31:0] pe3_lane5_strm0 [0:4095];
  reg [31:0] pe3_lane5_strm0_tmp     ;
  reg [31:0] pe3_lane5_strm1 [0:4095];
  reg [31:0] pe3_lane5_strm1_tmp     ;
  reg [31:0] pe3_lane6_strm0 [0:4095];
  reg [31:0] pe3_lane6_strm0_tmp     ;
  reg [31:0] pe3_lane6_strm1 [0:4095];
  reg [31:0] pe3_lane6_strm1_tmp     ;
  reg [31:0] pe3_lane7_strm0 [0:4095];
  reg [31:0] pe3_lane7_strm0_tmp     ;
  reg [31:0] pe3_lane7_strm1 [0:4095];
  reg [31:0] pe3_lane7_strm1_tmp     ;
  reg [31:0] pe3_lane8_strm0 [0:4095];
  reg [31:0] pe3_lane8_strm0_tmp     ;
  reg [31:0] pe3_lane8_strm1 [0:4095];
  reg [31:0] pe3_lane8_strm1_tmp     ;
  reg [31:0] pe3_lane9_strm0 [0:4095];
  reg [31:0] pe3_lane9_strm0_tmp     ;
  reg [31:0] pe3_lane9_strm1 [0:4095];
  reg [31:0] pe3_lane9_strm1_tmp     ;
  reg [31:0] pe3_lane10_strm0 [0:4095];
  reg [31:0] pe3_lane10_strm0_tmp     ;
  reg [31:0] pe3_lane10_strm1 [0:4095];
  reg [31:0] pe3_lane10_strm1_tmp     ;
  reg [31:0] pe3_lane11_strm0 [0:4095];
  reg [31:0] pe3_lane11_strm0_tmp     ;
  reg [31:0] pe3_lane11_strm1 [0:4095];
  reg [31:0] pe3_lane11_strm1_tmp     ;
  reg [31:0] pe3_lane12_strm0 [0:4095];
  reg [31:0] pe3_lane12_strm0_tmp     ;
  reg [31:0] pe3_lane12_strm1 [0:4095];
  reg [31:0] pe3_lane12_strm1_tmp     ;
  reg [31:0] pe3_lane13_strm0 [0:4095];
  reg [31:0] pe3_lane13_strm0_tmp     ;
  reg [31:0] pe3_lane13_strm1 [0:4095];
  reg [31:0] pe3_lane13_strm1_tmp     ;
  reg [31:0] pe3_lane14_strm0 [0:4095];
  reg [31:0] pe3_lane14_strm0_tmp     ;
  reg [31:0] pe3_lane14_strm1 [0:4095];
  reg [31:0] pe3_lane14_strm1_tmp     ;
  reg [31:0] pe3_lane15_strm0 [0:4095];
  reg [31:0] pe3_lane15_strm0_tmp     ;
  reg [31:0] pe3_lane15_strm1 [0:4095];
  reg [31:0] pe3_lane15_strm1_tmp     ;
  reg [31:0] pe3_lane16_strm0 [0:4095];
  reg [31:0] pe3_lane16_strm0_tmp     ;
  reg [31:0] pe3_lane16_strm1 [0:4095];
  reg [31:0] pe3_lane16_strm1_tmp     ;
  reg [31:0] pe3_lane17_strm0 [0:4095];
  reg [31:0] pe3_lane17_strm0_tmp     ;
  reg [31:0] pe3_lane17_strm1 [0:4095];
  reg [31:0] pe3_lane17_strm1_tmp     ;
  reg [31:0] pe3_lane18_strm0 [0:4095];
  reg [31:0] pe3_lane18_strm0_tmp     ;
  reg [31:0] pe3_lane18_strm1 [0:4095];
  reg [31:0] pe3_lane18_strm1_tmp     ;
  reg [31:0] pe3_lane19_strm0 [0:4095];
  reg [31:0] pe3_lane19_strm0_tmp     ;
  reg [31:0] pe3_lane19_strm1 [0:4095];
  reg [31:0] pe3_lane19_strm1_tmp     ;
  reg [31:0] pe3_lane20_strm0 [0:4095];
  reg [31:0] pe3_lane20_strm0_tmp     ;
  reg [31:0] pe3_lane20_strm1 [0:4095];
  reg [31:0] pe3_lane20_strm1_tmp     ;
  reg [31:0] pe3_lane21_strm0 [0:4095];
  reg [31:0] pe3_lane21_strm0_tmp     ;
  reg [31:0] pe3_lane21_strm1 [0:4095];
  reg [31:0] pe3_lane21_strm1_tmp     ;
  reg [31:0] pe3_lane22_strm0 [0:4095];
  reg [31:0] pe3_lane22_strm0_tmp     ;
  reg [31:0] pe3_lane22_strm1 [0:4095];
  reg [31:0] pe3_lane22_strm1_tmp     ;
  reg [31:0] pe3_lane23_strm0 [0:4095];
  reg [31:0] pe3_lane23_strm0_tmp     ;
  reg [31:0] pe3_lane23_strm1 [0:4095];
  reg [31:0] pe3_lane23_strm1_tmp     ;
  reg [31:0] pe3_lane24_strm0 [0:4095];
  reg [31:0] pe3_lane24_strm0_tmp     ;
  reg [31:0] pe3_lane24_strm1 [0:4095];
  reg [31:0] pe3_lane24_strm1_tmp     ;
  reg [31:0] pe3_lane25_strm0 [0:4095];
  reg [31:0] pe3_lane25_strm0_tmp     ;
  reg [31:0] pe3_lane25_strm1 [0:4095];
  reg [31:0] pe3_lane25_strm1_tmp     ;
  reg [31:0] pe3_lane26_strm0 [0:4095];
  reg [31:0] pe3_lane26_strm0_tmp     ;
  reg [31:0] pe3_lane26_strm1 [0:4095];
  reg [31:0] pe3_lane26_strm1_tmp     ;
  reg [31:0] pe3_lane27_strm0 [0:4095];
  reg [31:0] pe3_lane27_strm0_tmp     ;
  reg [31:0] pe3_lane27_strm1 [0:4095];
  reg [31:0] pe3_lane27_strm1_tmp     ;
  reg [31:0] pe3_lane28_strm0 [0:4095];
  reg [31:0] pe3_lane28_strm0_tmp     ;
  reg [31:0] pe3_lane28_strm1 [0:4095];
  reg [31:0] pe3_lane28_strm1_tmp     ;
  reg [31:0] pe3_lane29_strm0 [0:4095];
  reg [31:0] pe3_lane29_strm0_tmp     ;
  reg [31:0] pe3_lane29_strm1 [0:4095];
  reg [31:0] pe3_lane29_strm1_tmp     ;
  reg [31:0] pe3_lane30_strm0 [0:4095];
  reg [31:0] pe3_lane30_strm0_tmp     ;
  reg [31:0] pe3_lane30_strm1 [0:4095];
  reg [31:0] pe3_lane30_strm1_tmp     ;
  reg [31:0] pe3_lane31_strm0 [0:4095];
  reg [31:0] pe3_lane31_strm0_tmp     ;
  reg [31:0] pe3_lane31_strm1 [0:4095];
  reg [31:0] pe3_lane31_strm1_tmp     ;
  reg [31:0] pe4_lane0_strm0 [0:4095];
  reg [31:0] pe4_lane0_strm0_tmp     ;
  reg [31:0] pe4_lane0_strm1 [0:4095];
  reg [31:0] pe4_lane0_strm1_tmp     ;
  reg [31:0] pe4_lane1_strm0 [0:4095];
  reg [31:0] pe4_lane1_strm0_tmp     ;
  reg [31:0] pe4_lane1_strm1 [0:4095];
  reg [31:0] pe4_lane1_strm1_tmp     ;
  reg [31:0] pe4_lane2_strm0 [0:4095];
  reg [31:0] pe4_lane2_strm0_tmp     ;
  reg [31:0] pe4_lane2_strm1 [0:4095];
  reg [31:0] pe4_lane2_strm1_tmp     ;
  reg [31:0] pe4_lane3_strm0 [0:4095];
  reg [31:0] pe4_lane3_strm0_tmp     ;
  reg [31:0] pe4_lane3_strm1 [0:4095];
  reg [31:0] pe4_lane3_strm1_tmp     ;
  reg [31:0] pe4_lane4_strm0 [0:4095];
  reg [31:0] pe4_lane4_strm0_tmp     ;
  reg [31:0] pe4_lane4_strm1 [0:4095];
  reg [31:0] pe4_lane4_strm1_tmp     ;
  reg [31:0] pe4_lane5_strm0 [0:4095];
  reg [31:0] pe4_lane5_strm0_tmp     ;
  reg [31:0] pe4_lane5_strm1 [0:4095];
  reg [31:0] pe4_lane5_strm1_tmp     ;
  reg [31:0] pe4_lane6_strm0 [0:4095];
  reg [31:0] pe4_lane6_strm0_tmp     ;
  reg [31:0] pe4_lane6_strm1 [0:4095];
  reg [31:0] pe4_lane6_strm1_tmp     ;
  reg [31:0] pe4_lane7_strm0 [0:4095];
  reg [31:0] pe4_lane7_strm0_tmp     ;
  reg [31:0] pe4_lane7_strm1 [0:4095];
  reg [31:0] pe4_lane7_strm1_tmp     ;
  reg [31:0] pe4_lane8_strm0 [0:4095];
  reg [31:0] pe4_lane8_strm0_tmp     ;
  reg [31:0] pe4_lane8_strm1 [0:4095];
  reg [31:0] pe4_lane8_strm1_tmp     ;
  reg [31:0] pe4_lane9_strm0 [0:4095];
  reg [31:0] pe4_lane9_strm0_tmp     ;
  reg [31:0] pe4_lane9_strm1 [0:4095];
  reg [31:0] pe4_lane9_strm1_tmp     ;
  reg [31:0] pe4_lane10_strm0 [0:4095];
  reg [31:0] pe4_lane10_strm0_tmp     ;
  reg [31:0] pe4_lane10_strm1 [0:4095];
  reg [31:0] pe4_lane10_strm1_tmp     ;
  reg [31:0] pe4_lane11_strm0 [0:4095];
  reg [31:0] pe4_lane11_strm0_tmp     ;
  reg [31:0] pe4_lane11_strm1 [0:4095];
  reg [31:0] pe4_lane11_strm1_tmp     ;
  reg [31:0] pe4_lane12_strm0 [0:4095];
  reg [31:0] pe4_lane12_strm0_tmp     ;
  reg [31:0] pe4_lane12_strm1 [0:4095];
  reg [31:0] pe4_lane12_strm1_tmp     ;
  reg [31:0] pe4_lane13_strm0 [0:4095];
  reg [31:0] pe4_lane13_strm0_tmp     ;
  reg [31:0] pe4_lane13_strm1 [0:4095];
  reg [31:0] pe4_lane13_strm1_tmp     ;
  reg [31:0] pe4_lane14_strm0 [0:4095];
  reg [31:0] pe4_lane14_strm0_tmp     ;
  reg [31:0] pe4_lane14_strm1 [0:4095];
  reg [31:0] pe4_lane14_strm1_tmp     ;
  reg [31:0] pe4_lane15_strm0 [0:4095];
  reg [31:0] pe4_lane15_strm0_tmp     ;
  reg [31:0] pe4_lane15_strm1 [0:4095];
  reg [31:0] pe4_lane15_strm1_tmp     ;
  reg [31:0] pe4_lane16_strm0 [0:4095];
  reg [31:0] pe4_lane16_strm0_tmp     ;
  reg [31:0] pe4_lane16_strm1 [0:4095];
  reg [31:0] pe4_lane16_strm1_tmp     ;
  reg [31:0] pe4_lane17_strm0 [0:4095];
  reg [31:0] pe4_lane17_strm0_tmp     ;
  reg [31:0] pe4_lane17_strm1 [0:4095];
  reg [31:0] pe4_lane17_strm1_tmp     ;
  reg [31:0] pe4_lane18_strm0 [0:4095];
  reg [31:0] pe4_lane18_strm0_tmp     ;
  reg [31:0] pe4_lane18_strm1 [0:4095];
  reg [31:0] pe4_lane18_strm1_tmp     ;
  reg [31:0] pe4_lane19_strm0 [0:4095];
  reg [31:0] pe4_lane19_strm0_tmp     ;
  reg [31:0] pe4_lane19_strm1 [0:4095];
  reg [31:0] pe4_lane19_strm1_tmp     ;
  reg [31:0] pe4_lane20_strm0 [0:4095];
  reg [31:0] pe4_lane20_strm0_tmp     ;
  reg [31:0] pe4_lane20_strm1 [0:4095];
  reg [31:0] pe4_lane20_strm1_tmp     ;
  reg [31:0] pe4_lane21_strm0 [0:4095];
  reg [31:0] pe4_lane21_strm0_tmp     ;
  reg [31:0] pe4_lane21_strm1 [0:4095];
  reg [31:0] pe4_lane21_strm1_tmp     ;
  reg [31:0] pe4_lane22_strm0 [0:4095];
  reg [31:0] pe4_lane22_strm0_tmp     ;
  reg [31:0] pe4_lane22_strm1 [0:4095];
  reg [31:0] pe4_lane22_strm1_tmp     ;
  reg [31:0] pe4_lane23_strm0 [0:4095];
  reg [31:0] pe4_lane23_strm0_tmp     ;
  reg [31:0] pe4_lane23_strm1 [0:4095];
  reg [31:0] pe4_lane23_strm1_tmp     ;
  reg [31:0] pe4_lane24_strm0 [0:4095];
  reg [31:0] pe4_lane24_strm0_tmp     ;
  reg [31:0] pe4_lane24_strm1 [0:4095];
  reg [31:0] pe4_lane24_strm1_tmp     ;
  reg [31:0] pe4_lane25_strm0 [0:4095];
  reg [31:0] pe4_lane25_strm0_tmp     ;
  reg [31:0] pe4_lane25_strm1 [0:4095];
  reg [31:0] pe4_lane25_strm1_tmp     ;
  reg [31:0] pe4_lane26_strm0 [0:4095];
  reg [31:0] pe4_lane26_strm0_tmp     ;
  reg [31:0] pe4_lane26_strm1 [0:4095];
  reg [31:0] pe4_lane26_strm1_tmp     ;
  reg [31:0] pe4_lane27_strm0 [0:4095];
  reg [31:0] pe4_lane27_strm0_tmp     ;
  reg [31:0] pe4_lane27_strm1 [0:4095];
  reg [31:0] pe4_lane27_strm1_tmp     ;
  reg [31:0] pe4_lane28_strm0 [0:4095];
  reg [31:0] pe4_lane28_strm0_tmp     ;
  reg [31:0] pe4_lane28_strm1 [0:4095];
  reg [31:0] pe4_lane28_strm1_tmp     ;
  reg [31:0] pe4_lane29_strm0 [0:4095];
  reg [31:0] pe4_lane29_strm0_tmp     ;
  reg [31:0] pe4_lane29_strm1 [0:4095];
  reg [31:0] pe4_lane29_strm1_tmp     ;
  reg [31:0] pe4_lane30_strm0 [0:4095];
  reg [31:0] pe4_lane30_strm0_tmp     ;
  reg [31:0] pe4_lane30_strm1 [0:4095];
  reg [31:0] pe4_lane30_strm1_tmp     ;
  reg [31:0] pe4_lane31_strm0 [0:4095];
  reg [31:0] pe4_lane31_strm0_tmp     ;
  reg [31:0] pe4_lane31_strm1 [0:4095];
  reg [31:0] pe4_lane31_strm1_tmp     ;
  reg [31:0] pe5_lane0_strm0 [0:4095];
  reg [31:0] pe5_lane0_strm0_tmp     ;
  reg [31:0] pe5_lane0_strm1 [0:4095];
  reg [31:0] pe5_lane0_strm1_tmp     ;
  reg [31:0] pe5_lane1_strm0 [0:4095];
  reg [31:0] pe5_lane1_strm0_tmp     ;
  reg [31:0] pe5_lane1_strm1 [0:4095];
  reg [31:0] pe5_lane1_strm1_tmp     ;
  reg [31:0] pe5_lane2_strm0 [0:4095];
  reg [31:0] pe5_lane2_strm0_tmp     ;
  reg [31:0] pe5_lane2_strm1 [0:4095];
  reg [31:0] pe5_lane2_strm1_tmp     ;
  reg [31:0] pe5_lane3_strm0 [0:4095];
  reg [31:0] pe5_lane3_strm0_tmp     ;
  reg [31:0] pe5_lane3_strm1 [0:4095];
  reg [31:0] pe5_lane3_strm1_tmp     ;
  reg [31:0] pe5_lane4_strm0 [0:4095];
  reg [31:0] pe5_lane4_strm0_tmp     ;
  reg [31:0] pe5_lane4_strm1 [0:4095];
  reg [31:0] pe5_lane4_strm1_tmp     ;
  reg [31:0] pe5_lane5_strm0 [0:4095];
  reg [31:0] pe5_lane5_strm0_tmp     ;
  reg [31:0] pe5_lane5_strm1 [0:4095];
  reg [31:0] pe5_lane5_strm1_tmp     ;
  reg [31:0] pe5_lane6_strm0 [0:4095];
  reg [31:0] pe5_lane6_strm0_tmp     ;
  reg [31:0] pe5_lane6_strm1 [0:4095];
  reg [31:0] pe5_lane6_strm1_tmp     ;
  reg [31:0] pe5_lane7_strm0 [0:4095];
  reg [31:0] pe5_lane7_strm0_tmp     ;
  reg [31:0] pe5_lane7_strm1 [0:4095];
  reg [31:0] pe5_lane7_strm1_tmp     ;
  reg [31:0] pe5_lane8_strm0 [0:4095];
  reg [31:0] pe5_lane8_strm0_tmp     ;
  reg [31:0] pe5_lane8_strm1 [0:4095];
  reg [31:0] pe5_lane8_strm1_tmp     ;
  reg [31:0] pe5_lane9_strm0 [0:4095];
  reg [31:0] pe5_lane9_strm0_tmp     ;
  reg [31:0] pe5_lane9_strm1 [0:4095];
  reg [31:0] pe5_lane9_strm1_tmp     ;
  reg [31:0] pe5_lane10_strm0 [0:4095];
  reg [31:0] pe5_lane10_strm0_tmp     ;
  reg [31:0] pe5_lane10_strm1 [0:4095];
  reg [31:0] pe5_lane10_strm1_tmp     ;
  reg [31:0] pe5_lane11_strm0 [0:4095];
  reg [31:0] pe5_lane11_strm0_tmp     ;
  reg [31:0] pe5_lane11_strm1 [0:4095];
  reg [31:0] pe5_lane11_strm1_tmp     ;
  reg [31:0] pe5_lane12_strm0 [0:4095];
  reg [31:0] pe5_lane12_strm0_tmp     ;
  reg [31:0] pe5_lane12_strm1 [0:4095];
  reg [31:0] pe5_lane12_strm1_tmp     ;
  reg [31:0] pe5_lane13_strm0 [0:4095];
  reg [31:0] pe5_lane13_strm0_tmp     ;
  reg [31:0] pe5_lane13_strm1 [0:4095];
  reg [31:0] pe5_lane13_strm1_tmp     ;
  reg [31:0] pe5_lane14_strm0 [0:4095];
  reg [31:0] pe5_lane14_strm0_tmp     ;
  reg [31:0] pe5_lane14_strm1 [0:4095];
  reg [31:0] pe5_lane14_strm1_tmp     ;
  reg [31:0] pe5_lane15_strm0 [0:4095];
  reg [31:0] pe5_lane15_strm0_tmp     ;
  reg [31:0] pe5_lane15_strm1 [0:4095];
  reg [31:0] pe5_lane15_strm1_tmp     ;
  reg [31:0] pe5_lane16_strm0 [0:4095];
  reg [31:0] pe5_lane16_strm0_tmp     ;
  reg [31:0] pe5_lane16_strm1 [0:4095];
  reg [31:0] pe5_lane16_strm1_tmp     ;
  reg [31:0] pe5_lane17_strm0 [0:4095];
  reg [31:0] pe5_lane17_strm0_tmp     ;
  reg [31:0] pe5_lane17_strm1 [0:4095];
  reg [31:0] pe5_lane17_strm1_tmp     ;
  reg [31:0] pe5_lane18_strm0 [0:4095];
  reg [31:0] pe5_lane18_strm0_tmp     ;
  reg [31:0] pe5_lane18_strm1 [0:4095];
  reg [31:0] pe5_lane18_strm1_tmp     ;
  reg [31:0] pe5_lane19_strm0 [0:4095];
  reg [31:0] pe5_lane19_strm0_tmp     ;
  reg [31:0] pe5_lane19_strm1 [0:4095];
  reg [31:0] pe5_lane19_strm1_tmp     ;
  reg [31:0] pe5_lane20_strm0 [0:4095];
  reg [31:0] pe5_lane20_strm0_tmp     ;
  reg [31:0] pe5_lane20_strm1 [0:4095];
  reg [31:0] pe5_lane20_strm1_tmp     ;
  reg [31:0] pe5_lane21_strm0 [0:4095];
  reg [31:0] pe5_lane21_strm0_tmp     ;
  reg [31:0] pe5_lane21_strm1 [0:4095];
  reg [31:0] pe5_lane21_strm1_tmp     ;
  reg [31:0] pe5_lane22_strm0 [0:4095];
  reg [31:0] pe5_lane22_strm0_tmp     ;
  reg [31:0] pe5_lane22_strm1 [0:4095];
  reg [31:0] pe5_lane22_strm1_tmp     ;
  reg [31:0] pe5_lane23_strm0 [0:4095];
  reg [31:0] pe5_lane23_strm0_tmp     ;
  reg [31:0] pe5_lane23_strm1 [0:4095];
  reg [31:0] pe5_lane23_strm1_tmp     ;
  reg [31:0] pe5_lane24_strm0 [0:4095];
  reg [31:0] pe5_lane24_strm0_tmp     ;
  reg [31:0] pe5_lane24_strm1 [0:4095];
  reg [31:0] pe5_lane24_strm1_tmp     ;
  reg [31:0] pe5_lane25_strm0 [0:4095];
  reg [31:0] pe5_lane25_strm0_tmp     ;
  reg [31:0] pe5_lane25_strm1 [0:4095];
  reg [31:0] pe5_lane25_strm1_tmp     ;
  reg [31:0] pe5_lane26_strm0 [0:4095];
  reg [31:0] pe5_lane26_strm0_tmp     ;
  reg [31:0] pe5_lane26_strm1 [0:4095];
  reg [31:0] pe5_lane26_strm1_tmp     ;
  reg [31:0] pe5_lane27_strm0 [0:4095];
  reg [31:0] pe5_lane27_strm0_tmp     ;
  reg [31:0] pe5_lane27_strm1 [0:4095];
  reg [31:0] pe5_lane27_strm1_tmp     ;
  reg [31:0] pe5_lane28_strm0 [0:4095];
  reg [31:0] pe5_lane28_strm0_tmp     ;
  reg [31:0] pe5_lane28_strm1 [0:4095];
  reg [31:0] pe5_lane28_strm1_tmp     ;
  reg [31:0] pe5_lane29_strm0 [0:4095];
  reg [31:0] pe5_lane29_strm0_tmp     ;
  reg [31:0] pe5_lane29_strm1 [0:4095];
  reg [31:0] pe5_lane29_strm1_tmp     ;
  reg [31:0] pe5_lane30_strm0 [0:4095];
  reg [31:0] pe5_lane30_strm0_tmp     ;
  reg [31:0] pe5_lane30_strm1 [0:4095];
  reg [31:0] pe5_lane30_strm1_tmp     ;
  reg [31:0] pe5_lane31_strm0 [0:4095];
  reg [31:0] pe5_lane31_strm0_tmp     ;
  reg [31:0] pe5_lane31_strm1 [0:4095];
  reg [31:0] pe5_lane31_strm1_tmp     ;
  reg [31:0] pe6_lane0_strm0 [0:4095];
  reg [31:0] pe6_lane0_strm0_tmp     ;
  reg [31:0] pe6_lane0_strm1 [0:4095];
  reg [31:0] pe6_lane0_strm1_tmp     ;
  reg [31:0] pe6_lane1_strm0 [0:4095];
  reg [31:0] pe6_lane1_strm0_tmp     ;
  reg [31:0] pe6_lane1_strm1 [0:4095];
  reg [31:0] pe6_lane1_strm1_tmp     ;
  reg [31:0] pe6_lane2_strm0 [0:4095];
  reg [31:0] pe6_lane2_strm0_tmp     ;
  reg [31:0] pe6_lane2_strm1 [0:4095];
  reg [31:0] pe6_lane2_strm1_tmp     ;
  reg [31:0] pe6_lane3_strm0 [0:4095];
  reg [31:0] pe6_lane3_strm0_tmp     ;
  reg [31:0] pe6_lane3_strm1 [0:4095];
  reg [31:0] pe6_lane3_strm1_tmp     ;
  reg [31:0] pe6_lane4_strm0 [0:4095];
  reg [31:0] pe6_lane4_strm0_tmp     ;
  reg [31:0] pe6_lane4_strm1 [0:4095];
  reg [31:0] pe6_lane4_strm1_tmp     ;
  reg [31:0] pe6_lane5_strm0 [0:4095];
  reg [31:0] pe6_lane5_strm0_tmp     ;
  reg [31:0] pe6_lane5_strm1 [0:4095];
  reg [31:0] pe6_lane5_strm1_tmp     ;
  reg [31:0] pe6_lane6_strm0 [0:4095];
  reg [31:0] pe6_lane6_strm0_tmp     ;
  reg [31:0] pe6_lane6_strm1 [0:4095];
  reg [31:0] pe6_lane6_strm1_tmp     ;
  reg [31:0] pe6_lane7_strm0 [0:4095];
  reg [31:0] pe6_lane7_strm0_tmp     ;
  reg [31:0] pe6_lane7_strm1 [0:4095];
  reg [31:0] pe6_lane7_strm1_tmp     ;
  reg [31:0] pe6_lane8_strm0 [0:4095];
  reg [31:0] pe6_lane8_strm0_tmp     ;
  reg [31:0] pe6_lane8_strm1 [0:4095];
  reg [31:0] pe6_lane8_strm1_tmp     ;
  reg [31:0] pe6_lane9_strm0 [0:4095];
  reg [31:0] pe6_lane9_strm0_tmp     ;
  reg [31:0] pe6_lane9_strm1 [0:4095];
  reg [31:0] pe6_lane9_strm1_tmp     ;
  reg [31:0] pe6_lane10_strm0 [0:4095];
  reg [31:0] pe6_lane10_strm0_tmp     ;
  reg [31:0] pe6_lane10_strm1 [0:4095];
  reg [31:0] pe6_lane10_strm1_tmp     ;
  reg [31:0] pe6_lane11_strm0 [0:4095];
  reg [31:0] pe6_lane11_strm0_tmp     ;
  reg [31:0] pe6_lane11_strm1 [0:4095];
  reg [31:0] pe6_lane11_strm1_tmp     ;
  reg [31:0] pe6_lane12_strm0 [0:4095];
  reg [31:0] pe6_lane12_strm0_tmp     ;
  reg [31:0] pe6_lane12_strm1 [0:4095];
  reg [31:0] pe6_lane12_strm1_tmp     ;
  reg [31:0] pe6_lane13_strm0 [0:4095];
  reg [31:0] pe6_lane13_strm0_tmp     ;
  reg [31:0] pe6_lane13_strm1 [0:4095];
  reg [31:0] pe6_lane13_strm1_tmp     ;
  reg [31:0] pe6_lane14_strm0 [0:4095];
  reg [31:0] pe6_lane14_strm0_tmp     ;
  reg [31:0] pe6_lane14_strm1 [0:4095];
  reg [31:0] pe6_lane14_strm1_tmp     ;
  reg [31:0] pe6_lane15_strm0 [0:4095];
  reg [31:0] pe6_lane15_strm0_tmp     ;
  reg [31:0] pe6_lane15_strm1 [0:4095];
  reg [31:0] pe6_lane15_strm1_tmp     ;
  reg [31:0] pe6_lane16_strm0 [0:4095];
  reg [31:0] pe6_lane16_strm0_tmp     ;
  reg [31:0] pe6_lane16_strm1 [0:4095];
  reg [31:0] pe6_lane16_strm1_tmp     ;
  reg [31:0] pe6_lane17_strm0 [0:4095];
  reg [31:0] pe6_lane17_strm0_tmp     ;
  reg [31:0] pe6_lane17_strm1 [0:4095];
  reg [31:0] pe6_lane17_strm1_tmp     ;
  reg [31:0] pe6_lane18_strm0 [0:4095];
  reg [31:0] pe6_lane18_strm0_tmp     ;
  reg [31:0] pe6_lane18_strm1 [0:4095];
  reg [31:0] pe6_lane18_strm1_tmp     ;
  reg [31:0] pe6_lane19_strm0 [0:4095];
  reg [31:0] pe6_lane19_strm0_tmp     ;
  reg [31:0] pe6_lane19_strm1 [0:4095];
  reg [31:0] pe6_lane19_strm1_tmp     ;
  reg [31:0] pe6_lane20_strm0 [0:4095];
  reg [31:0] pe6_lane20_strm0_tmp     ;
  reg [31:0] pe6_lane20_strm1 [0:4095];
  reg [31:0] pe6_lane20_strm1_tmp     ;
  reg [31:0] pe6_lane21_strm0 [0:4095];
  reg [31:0] pe6_lane21_strm0_tmp     ;
  reg [31:0] pe6_lane21_strm1 [0:4095];
  reg [31:0] pe6_lane21_strm1_tmp     ;
  reg [31:0] pe6_lane22_strm0 [0:4095];
  reg [31:0] pe6_lane22_strm0_tmp     ;
  reg [31:0] pe6_lane22_strm1 [0:4095];
  reg [31:0] pe6_lane22_strm1_tmp     ;
  reg [31:0] pe6_lane23_strm0 [0:4095];
  reg [31:0] pe6_lane23_strm0_tmp     ;
  reg [31:0] pe6_lane23_strm1 [0:4095];
  reg [31:0] pe6_lane23_strm1_tmp     ;
  reg [31:0] pe6_lane24_strm0 [0:4095];
  reg [31:0] pe6_lane24_strm0_tmp     ;
  reg [31:0] pe6_lane24_strm1 [0:4095];
  reg [31:0] pe6_lane24_strm1_tmp     ;
  reg [31:0] pe6_lane25_strm0 [0:4095];
  reg [31:0] pe6_lane25_strm0_tmp     ;
  reg [31:0] pe6_lane25_strm1 [0:4095];
  reg [31:0] pe6_lane25_strm1_tmp     ;
  reg [31:0] pe6_lane26_strm0 [0:4095];
  reg [31:0] pe6_lane26_strm0_tmp     ;
  reg [31:0] pe6_lane26_strm1 [0:4095];
  reg [31:0] pe6_lane26_strm1_tmp     ;
  reg [31:0] pe6_lane27_strm0 [0:4095];
  reg [31:0] pe6_lane27_strm0_tmp     ;
  reg [31:0] pe6_lane27_strm1 [0:4095];
  reg [31:0] pe6_lane27_strm1_tmp     ;
  reg [31:0] pe6_lane28_strm0 [0:4095];
  reg [31:0] pe6_lane28_strm0_tmp     ;
  reg [31:0] pe6_lane28_strm1 [0:4095];
  reg [31:0] pe6_lane28_strm1_tmp     ;
  reg [31:0] pe6_lane29_strm0 [0:4095];
  reg [31:0] pe6_lane29_strm0_tmp     ;
  reg [31:0] pe6_lane29_strm1 [0:4095];
  reg [31:0] pe6_lane29_strm1_tmp     ;
  reg [31:0] pe6_lane30_strm0 [0:4095];
  reg [31:0] pe6_lane30_strm0_tmp     ;
  reg [31:0] pe6_lane30_strm1 [0:4095];
  reg [31:0] pe6_lane30_strm1_tmp     ;
  reg [31:0] pe6_lane31_strm0 [0:4095];
  reg [31:0] pe6_lane31_strm0_tmp     ;
  reg [31:0] pe6_lane31_strm1 [0:4095];
  reg [31:0] pe6_lane31_strm1_tmp     ;
  reg [31:0] pe7_lane0_strm0 [0:4095];
  reg [31:0] pe7_lane0_strm0_tmp     ;
  reg [31:0] pe7_lane0_strm1 [0:4095];
  reg [31:0] pe7_lane0_strm1_tmp     ;
  reg [31:0] pe7_lane1_strm0 [0:4095];
  reg [31:0] pe7_lane1_strm0_tmp     ;
  reg [31:0] pe7_lane1_strm1 [0:4095];
  reg [31:0] pe7_lane1_strm1_tmp     ;
  reg [31:0] pe7_lane2_strm0 [0:4095];
  reg [31:0] pe7_lane2_strm0_tmp     ;
  reg [31:0] pe7_lane2_strm1 [0:4095];
  reg [31:0] pe7_lane2_strm1_tmp     ;
  reg [31:0] pe7_lane3_strm0 [0:4095];
  reg [31:0] pe7_lane3_strm0_tmp     ;
  reg [31:0] pe7_lane3_strm1 [0:4095];
  reg [31:0] pe7_lane3_strm1_tmp     ;
  reg [31:0] pe7_lane4_strm0 [0:4095];
  reg [31:0] pe7_lane4_strm0_tmp     ;
  reg [31:0] pe7_lane4_strm1 [0:4095];
  reg [31:0] pe7_lane4_strm1_tmp     ;
  reg [31:0] pe7_lane5_strm0 [0:4095];
  reg [31:0] pe7_lane5_strm0_tmp     ;
  reg [31:0] pe7_lane5_strm1 [0:4095];
  reg [31:0] pe7_lane5_strm1_tmp     ;
  reg [31:0] pe7_lane6_strm0 [0:4095];
  reg [31:0] pe7_lane6_strm0_tmp     ;
  reg [31:0] pe7_lane6_strm1 [0:4095];
  reg [31:0] pe7_lane6_strm1_tmp     ;
  reg [31:0] pe7_lane7_strm0 [0:4095];
  reg [31:0] pe7_lane7_strm0_tmp     ;
  reg [31:0] pe7_lane7_strm1 [0:4095];
  reg [31:0] pe7_lane7_strm1_tmp     ;
  reg [31:0] pe7_lane8_strm0 [0:4095];
  reg [31:0] pe7_lane8_strm0_tmp     ;
  reg [31:0] pe7_lane8_strm1 [0:4095];
  reg [31:0] pe7_lane8_strm1_tmp     ;
  reg [31:0] pe7_lane9_strm0 [0:4095];
  reg [31:0] pe7_lane9_strm0_tmp     ;
  reg [31:0] pe7_lane9_strm1 [0:4095];
  reg [31:0] pe7_lane9_strm1_tmp     ;
  reg [31:0] pe7_lane10_strm0 [0:4095];
  reg [31:0] pe7_lane10_strm0_tmp     ;
  reg [31:0] pe7_lane10_strm1 [0:4095];
  reg [31:0] pe7_lane10_strm1_tmp     ;
  reg [31:0] pe7_lane11_strm0 [0:4095];
  reg [31:0] pe7_lane11_strm0_tmp     ;
  reg [31:0] pe7_lane11_strm1 [0:4095];
  reg [31:0] pe7_lane11_strm1_tmp     ;
  reg [31:0] pe7_lane12_strm0 [0:4095];
  reg [31:0] pe7_lane12_strm0_tmp     ;
  reg [31:0] pe7_lane12_strm1 [0:4095];
  reg [31:0] pe7_lane12_strm1_tmp     ;
  reg [31:0] pe7_lane13_strm0 [0:4095];
  reg [31:0] pe7_lane13_strm0_tmp     ;
  reg [31:0] pe7_lane13_strm1 [0:4095];
  reg [31:0] pe7_lane13_strm1_tmp     ;
  reg [31:0] pe7_lane14_strm0 [0:4095];
  reg [31:0] pe7_lane14_strm0_tmp     ;
  reg [31:0] pe7_lane14_strm1 [0:4095];
  reg [31:0] pe7_lane14_strm1_tmp     ;
  reg [31:0] pe7_lane15_strm0 [0:4095];
  reg [31:0] pe7_lane15_strm0_tmp     ;
  reg [31:0] pe7_lane15_strm1 [0:4095];
  reg [31:0] pe7_lane15_strm1_tmp     ;
  reg [31:0] pe7_lane16_strm0 [0:4095];
  reg [31:0] pe7_lane16_strm0_tmp     ;
  reg [31:0] pe7_lane16_strm1 [0:4095];
  reg [31:0] pe7_lane16_strm1_tmp     ;
  reg [31:0] pe7_lane17_strm0 [0:4095];
  reg [31:0] pe7_lane17_strm0_tmp     ;
  reg [31:0] pe7_lane17_strm1 [0:4095];
  reg [31:0] pe7_lane17_strm1_tmp     ;
  reg [31:0] pe7_lane18_strm0 [0:4095];
  reg [31:0] pe7_lane18_strm0_tmp     ;
  reg [31:0] pe7_lane18_strm1 [0:4095];
  reg [31:0] pe7_lane18_strm1_tmp     ;
  reg [31:0] pe7_lane19_strm0 [0:4095];
  reg [31:0] pe7_lane19_strm0_tmp     ;
  reg [31:0] pe7_lane19_strm1 [0:4095];
  reg [31:0] pe7_lane19_strm1_tmp     ;
  reg [31:0] pe7_lane20_strm0 [0:4095];
  reg [31:0] pe7_lane20_strm0_tmp     ;
  reg [31:0] pe7_lane20_strm1 [0:4095];
  reg [31:0] pe7_lane20_strm1_tmp     ;
  reg [31:0] pe7_lane21_strm0 [0:4095];
  reg [31:0] pe7_lane21_strm0_tmp     ;
  reg [31:0] pe7_lane21_strm1 [0:4095];
  reg [31:0] pe7_lane21_strm1_tmp     ;
  reg [31:0] pe7_lane22_strm0 [0:4095];
  reg [31:0] pe7_lane22_strm0_tmp     ;
  reg [31:0] pe7_lane22_strm1 [0:4095];
  reg [31:0] pe7_lane22_strm1_tmp     ;
  reg [31:0] pe7_lane23_strm0 [0:4095];
  reg [31:0] pe7_lane23_strm0_tmp     ;
  reg [31:0] pe7_lane23_strm1 [0:4095];
  reg [31:0] pe7_lane23_strm1_tmp     ;
  reg [31:0] pe7_lane24_strm0 [0:4095];
  reg [31:0] pe7_lane24_strm0_tmp     ;
  reg [31:0] pe7_lane24_strm1 [0:4095];
  reg [31:0] pe7_lane24_strm1_tmp     ;
  reg [31:0] pe7_lane25_strm0 [0:4095];
  reg [31:0] pe7_lane25_strm0_tmp     ;
  reg [31:0] pe7_lane25_strm1 [0:4095];
  reg [31:0] pe7_lane25_strm1_tmp     ;
  reg [31:0] pe7_lane26_strm0 [0:4095];
  reg [31:0] pe7_lane26_strm0_tmp     ;
  reg [31:0] pe7_lane26_strm1 [0:4095];
  reg [31:0] pe7_lane26_strm1_tmp     ;
  reg [31:0] pe7_lane27_strm0 [0:4095];
  reg [31:0] pe7_lane27_strm0_tmp     ;
  reg [31:0] pe7_lane27_strm1 [0:4095];
  reg [31:0] pe7_lane27_strm1_tmp     ;
  reg [31:0] pe7_lane28_strm0 [0:4095];
  reg [31:0] pe7_lane28_strm0_tmp     ;
  reg [31:0] pe7_lane28_strm1 [0:4095];
  reg [31:0] pe7_lane28_strm1_tmp     ;
  reg [31:0] pe7_lane29_strm0 [0:4095];
  reg [31:0] pe7_lane29_strm0_tmp     ;
  reg [31:0] pe7_lane29_strm1 [0:4095];
  reg [31:0] pe7_lane29_strm1_tmp     ;
  reg [31:0] pe7_lane30_strm0 [0:4095];
  reg [31:0] pe7_lane30_strm0_tmp     ;
  reg [31:0] pe7_lane30_strm1 [0:4095];
  reg [31:0] pe7_lane30_strm1_tmp     ;
  reg [31:0] pe7_lane31_strm0 [0:4095];
  reg [31:0] pe7_lane31_strm0_tmp     ;
  reg [31:0] pe7_lane31_strm1 [0:4095];
  reg [31:0] pe7_lane31_strm1_tmp     ;
  reg [31:0] pe8_lane0_strm0 [0:4095];
  reg [31:0] pe8_lane0_strm0_tmp     ;
  reg [31:0] pe8_lane0_strm1 [0:4095];
  reg [31:0] pe8_lane0_strm1_tmp     ;
  reg [31:0] pe8_lane1_strm0 [0:4095];
  reg [31:0] pe8_lane1_strm0_tmp     ;
  reg [31:0] pe8_lane1_strm1 [0:4095];
  reg [31:0] pe8_lane1_strm1_tmp     ;
  reg [31:0] pe8_lane2_strm0 [0:4095];
  reg [31:0] pe8_lane2_strm0_tmp     ;
  reg [31:0] pe8_lane2_strm1 [0:4095];
  reg [31:0] pe8_lane2_strm1_tmp     ;
  reg [31:0] pe8_lane3_strm0 [0:4095];
  reg [31:0] pe8_lane3_strm0_tmp     ;
  reg [31:0] pe8_lane3_strm1 [0:4095];
  reg [31:0] pe8_lane3_strm1_tmp     ;
  reg [31:0] pe8_lane4_strm0 [0:4095];
  reg [31:0] pe8_lane4_strm0_tmp     ;
  reg [31:0] pe8_lane4_strm1 [0:4095];
  reg [31:0] pe8_lane4_strm1_tmp     ;
  reg [31:0] pe8_lane5_strm0 [0:4095];
  reg [31:0] pe8_lane5_strm0_tmp     ;
  reg [31:0] pe8_lane5_strm1 [0:4095];
  reg [31:0] pe8_lane5_strm1_tmp     ;
  reg [31:0] pe8_lane6_strm0 [0:4095];
  reg [31:0] pe8_lane6_strm0_tmp     ;
  reg [31:0] pe8_lane6_strm1 [0:4095];
  reg [31:0] pe8_lane6_strm1_tmp     ;
  reg [31:0] pe8_lane7_strm0 [0:4095];
  reg [31:0] pe8_lane7_strm0_tmp     ;
  reg [31:0] pe8_lane7_strm1 [0:4095];
  reg [31:0] pe8_lane7_strm1_tmp     ;
  reg [31:0] pe8_lane8_strm0 [0:4095];
  reg [31:0] pe8_lane8_strm0_tmp     ;
  reg [31:0] pe8_lane8_strm1 [0:4095];
  reg [31:0] pe8_lane8_strm1_tmp     ;
  reg [31:0] pe8_lane9_strm0 [0:4095];
  reg [31:0] pe8_lane9_strm0_tmp     ;
  reg [31:0] pe8_lane9_strm1 [0:4095];
  reg [31:0] pe8_lane9_strm1_tmp     ;
  reg [31:0] pe8_lane10_strm0 [0:4095];
  reg [31:0] pe8_lane10_strm0_tmp     ;
  reg [31:0] pe8_lane10_strm1 [0:4095];
  reg [31:0] pe8_lane10_strm1_tmp     ;
  reg [31:0] pe8_lane11_strm0 [0:4095];
  reg [31:0] pe8_lane11_strm0_tmp     ;
  reg [31:0] pe8_lane11_strm1 [0:4095];
  reg [31:0] pe8_lane11_strm1_tmp     ;
  reg [31:0] pe8_lane12_strm0 [0:4095];
  reg [31:0] pe8_lane12_strm0_tmp     ;
  reg [31:0] pe8_lane12_strm1 [0:4095];
  reg [31:0] pe8_lane12_strm1_tmp     ;
  reg [31:0] pe8_lane13_strm0 [0:4095];
  reg [31:0] pe8_lane13_strm0_tmp     ;
  reg [31:0] pe8_lane13_strm1 [0:4095];
  reg [31:0] pe8_lane13_strm1_tmp     ;
  reg [31:0] pe8_lane14_strm0 [0:4095];
  reg [31:0] pe8_lane14_strm0_tmp     ;
  reg [31:0] pe8_lane14_strm1 [0:4095];
  reg [31:0] pe8_lane14_strm1_tmp     ;
  reg [31:0] pe8_lane15_strm0 [0:4095];
  reg [31:0] pe8_lane15_strm0_tmp     ;
  reg [31:0] pe8_lane15_strm1 [0:4095];
  reg [31:0] pe8_lane15_strm1_tmp     ;
  reg [31:0] pe8_lane16_strm0 [0:4095];
  reg [31:0] pe8_lane16_strm0_tmp     ;
  reg [31:0] pe8_lane16_strm1 [0:4095];
  reg [31:0] pe8_lane16_strm1_tmp     ;
  reg [31:0] pe8_lane17_strm0 [0:4095];
  reg [31:0] pe8_lane17_strm0_tmp     ;
  reg [31:0] pe8_lane17_strm1 [0:4095];
  reg [31:0] pe8_lane17_strm1_tmp     ;
  reg [31:0] pe8_lane18_strm0 [0:4095];
  reg [31:0] pe8_lane18_strm0_tmp     ;
  reg [31:0] pe8_lane18_strm1 [0:4095];
  reg [31:0] pe8_lane18_strm1_tmp     ;
  reg [31:0] pe8_lane19_strm0 [0:4095];
  reg [31:0] pe8_lane19_strm0_tmp     ;
  reg [31:0] pe8_lane19_strm1 [0:4095];
  reg [31:0] pe8_lane19_strm1_tmp     ;
  reg [31:0] pe8_lane20_strm0 [0:4095];
  reg [31:0] pe8_lane20_strm0_tmp     ;
  reg [31:0] pe8_lane20_strm1 [0:4095];
  reg [31:0] pe8_lane20_strm1_tmp     ;
  reg [31:0] pe8_lane21_strm0 [0:4095];
  reg [31:0] pe8_lane21_strm0_tmp     ;
  reg [31:0] pe8_lane21_strm1 [0:4095];
  reg [31:0] pe8_lane21_strm1_tmp     ;
  reg [31:0] pe8_lane22_strm0 [0:4095];
  reg [31:0] pe8_lane22_strm0_tmp     ;
  reg [31:0] pe8_lane22_strm1 [0:4095];
  reg [31:0] pe8_lane22_strm1_tmp     ;
  reg [31:0] pe8_lane23_strm0 [0:4095];
  reg [31:0] pe8_lane23_strm0_tmp     ;
  reg [31:0] pe8_lane23_strm1 [0:4095];
  reg [31:0] pe8_lane23_strm1_tmp     ;
  reg [31:0] pe8_lane24_strm0 [0:4095];
  reg [31:0] pe8_lane24_strm0_tmp     ;
  reg [31:0] pe8_lane24_strm1 [0:4095];
  reg [31:0] pe8_lane24_strm1_tmp     ;
  reg [31:0] pe8_lane25_strm0 [0:4095];
  reg [31:0] pe8_lane25_strm0_tmp     ;
  reg [31:0] pe8_lane25_strm1 [0:4095];
  reg [31:0] pe8_lane25_strm1_tmp     ;
  reg [31:0] pe8_lane26_strm0 [0:4095];
  reg [31:0] pe8_lane26_strm0_tmp     ;
  reg [31:0] pe8_lane26_strm1 [0:4095];
  reg [31:0] pe8_lane26_strm1_tmp     ;
  reg [31:0] pe8_lane27_strm0 [0:4095];
  reg [31:0] pe8_lane27_strm0_tmp     ;
  reg [31:0] pe8_lane27_strm1 [0:4095];
  reg [31:0] pe8_lane27_strm1_tmp     ;
  reg [31:0] pe8_lane28_strm0 [0:4095];
  reg [31:0] pe8_lane28_strm0_tmp     ;
  reg [31:0] pe8_lane28_strm1 [0:4095];
  reg [31:0] pe8_lane28_strm1_tmp     ;
  reg [31:0] pe8_lane29_strm0 [0:4095];
  reg [31:0] pe8_lane29_strm0_tmp     ;
  reg [31:0] pe8_lane29_strm1 [0:4095];
  reg [31:0] pe8_lane29_strm1_tmp     ;
  reg [31:0] pe8_lane30_strm0 [0:4095];
  reg [31:0] pe8_lane30_strm0_tmp     ;
  reg [31:0] pe8_lane30_strm1 [0:4095];
  reg [31:0] pe8_lane30_strm1_tmp     ;
  reg [31:0] pe8_lane31_strm0 [0:4095];
  reg [31:0] pe8_lane31_strm0_tmp     ;
  reg [31:0] pe8_lane31_strm1 [0:4095];
  reg [31:0] pe8_lane31_strm1_tmp     ;
  reg [31:0] pe9_lane0_strm0 [0:4095];
  reg [31:0] pe9_lane0_strm0_tmp     ;
  reg [31:0] pe9_lane0_strm1 [0:4095];
  reg [31:0] pe9_lane0_strm1_tmp     ;
  reg [31:0] pe9_lane1_strm0 [0:4095];
  reg [31:0] pe9_lane1_strm0_tmp     ;
  reg [31:0] pe9_lane1_strm1 [0:4095];
  reg [31:0] pe9_lane1_strm1_tmp     ;
  reg [31:0] pe9_lane2_strm0 [0:4095];
  reg [31:0] pe9_lane2_strm0_tmp     ;
  reg [31:0] pe9_lane2_strm1 [0:4095];
  reg [31:0] pe9_lane2_strm1_tmp     ;
  reg [31:0] pe9_lane3_strm0 [0:4095];
  reg [31:0] pe9_lane3_strm0_tmp     ;
  reg [31:0] pe9_lane3_strm1 [0:4095];
  reg [31:0] pe9_lane3_strm1_tmp     ;
  reg [31:0] pe9_lane4_strm0 [0:4095];
  reg [31:0] pe9_lane4_strm0_tmp     ;
  reg [31:0] pe9_lane4_strm1 [0:4095];
  reg [31:0] pe9_lane4_strm1_tmp     ;
  reg [31:0] pe9_lane5_strm0 [0:4095];
  reg [31:0] pe9_lane5_strm0_tmp     ;
  reg [31:0] pe9_lane5_strm1 [0:4095];
  reg [31:0] pe9_lane5_strm1_tmp     ;
  reg [31:0] pe9_lane6_strm0 [0:4095];
  reg [31:0] pe9_lane6_strm0_tmp     ;
  reg [31:0] pe9_lane6_strm1 [0:4095];
  reg [31:0] pe9_lane6_strm1_tmp     ;
  reg [31:0] pe9_lane7_strm0 [0:4095];
  reg [31:0] pe9_lane7_strm0_tmp     ;
  reg [31:0] pe9_lane7_strm1 [0:4095];
  reg [31:0] pe9_lane7_strm1_tmp     ;
  reg [31:0] pe9_lane8_strm0 [0:4095];
  reg [31:0] pe9_lane8_strm0_tmp     ;
  reg [31:0] pe9_lane8_strm1 [0:4095];
  reg [31:0] pe9_lane8_strm1_tmp     ;
  reg [31:0] pe9_lane9_strm0 [0:4095];
  reg [31:0] pe9_lane9_strm0_tmp     ;
  reg [31:0] pe9_lane9_strm1 [0:4095];
  reg [31:0] pe9_lane9_strm1_tmp     ;
  reg [31:0] pe9_lane10_strm0 [0:4095];
  reg [31:0] pe9_lane10_strm0_tmp     ;
  reg [31:0] pe9_lane10_strm1 [0:4095];
  reg [31:0] pe9_lane10_strm1_tmp     ;
  reg [31:0] pe9_lane11_strm0 [0:4095];
  reg [31:0] pe9_lane11_strm0_tmp     ;
  reg [31:0] pe9_lane11_strm1 [0:4095];
  reg [31:0] pe9_lane11_strm1_tmp     ;
  reg [31:0] pe9_lane12_strm0 [0:4095];
  reg [31:0] pe9_lane12_strm0_tmp     ;
  reg [31:0] pe9_lane12_strm1 [0:4095];
  reg [31:0] pe9_lane12_strm1_tmp     ;
  reg [31:0] pe9_lane13_strm0 [0:4095];
  reg [31:0] pe9_lane13_strm0_tmp     ;
  reg [31:0] pe9_lane13_strm1 [0:4095];
  reg [31:0] pe9_lane13_strm1_tmp     ;
  reg [31:0] pe9_lane14_strm0 [0:4095];
  reg [31:0] pe9_lane14_strm0_tmp     ;
  reg [31:0] pe9_lane14_strm1 [0:4095];
  reg [31:0] pe9_lane14_strm1_tmp     ;
  reg [31:0] pe9_lane15_strm0 [0:4095];
  reg [31:0] pe9_lane15_strm0_tmp     ;
  reg [31:0] pe9_lane15_strm1 [0:4095];
  reg [31:0] pe9_lane15_strm1_tmp     ;
  reg [31:0] pe9_lane16_strm0 [0:4095];
  reg [31:0] pe9_lane16_strm0_tmp     ;
  reg [31:0] pe9_lane16_strm1 [0:4095];
  reg [31:0] pe9_lane16_strm1_tmp     ;
  reg [31:0] pe9_lane17_strm0 [0:4095];
  reg [31:0] pe9_lane17_strm0_tmp     ;
  reg [31:0] pe9_lane17_strm1 [0:4095];
  reg [31:0] pe9_lane17_strm1_tmp     ;
  reg [31:0] pe9_lane18_strm0 [0:4095];
  reg [31:0] pe9_lane18_strm0_tmp     ;
  reg [31:0] pe9_lane18_strm1 [0:4095];
  reg [31:0] pe9_lane18_strm1_tmp     ;
  reg [31:0] pe9_lane19_strm0 [0:4095];
  reg [31:0] pe9_lane19_strm0_tmp     ;
  reg [31:0] pe9_lane19_strm1 [0:4095];
  reg [31:0] pe9_lane19_strm1_tmp     ;
  reg [31:0] pe9_lane20_strm0 [0:4095];
  reg [31:0] pe9_lane20_strm0_tmp     ;
  reg [31:0] pe9_lane20_strm1 [0:4095];
  reg [31:0] pe9_lane20_strm1_tmp     ;
  reg [31:0] pe9_lane21_strm0 [0:4095];
  reg [31:0] pe9_lane21_strm0_tmp     ;
  reg [31:0] pe9_lane21_strm1 [0:4095];
  reg [31:0] pe9_lane21_strm1_tmp     ;
  reg [31:0] pe9_lane22_strm0 [0:4095];
  reg [31:0] pe9_lane22_strm0_tmp     ;
  reg [31:0] pe9_lane22_strm1 [0:4095];
  reg [31:0] pe9_lane22_strm1_tmp     ;
  reg [31:0] pe9_lane23_strm0 [0:4095];
  reg [31:0] pe9_lane23_strm0_tmp     ;
  reg [31:0] pe9_lane23_strm1 [0:4095];
  reg [31:0] pe9_lane23_strm1_tmp     ;
  reg [31:0] pe9_lane24_strm0 [0:4095];
  reg [31:0] pe9_lane24_strm0_tmp     ;
  reg [31:0] pe9_lane24_strm1 [0:4095];
  reg [31:0] pe9_lane24_strm1_tmp     ;
  reg [31:0] pe9_lane25_strm0 [0:4095];
  reg [31:0] pe9_lane25_strm0_tmp     ;
  reg [31:0] pe9_lane25_strm1 [0:4095];
  reg [31:0] pe9_lane25_strm1_tmp     ;
  reg [31:0] pe9_lane26_strm0 [0:4095];
  reg [31:0] pe9_lane26_strm0_tmp     ;
  reg [31:0] pe9_lane26_strm1 [0:4095];
  reg [31:0] pe9_lane26_strm1_tmp     ;
  reg [31:0] pe9_lane27_strm0 [0:4095];
  reg [31:0] pe9_lane27_strm0_tmp     ;
  reg [31:0] pe9_lane27_strm1 [0:4095];
  reg [31:0] pe9_lane27_strm1_tmp     ;
  reg [31:0] pe9_lane28_strm0 [0:4095];
  reg [31:0] pe9_lane28_strm0_tmp     ;
  reg [31:0] pe9_lane28_strm1 [0:4095];
  reg [31:0] pe9_lane28_strm1_tmp     ;
  reg [31:0] pe9_lane29_strm0 [0:4095];
  reg [31:0] pe9_lane29_strm0_tmp     ;
  reg [31:0] pe9_lane29_strm1 [0:4095];
  reg [31:0] pe9_lane29_strm1_tmp     ;
  reg [31:0] pe9_lane30_strm0 [0:4095];
  reg [31:0] pe9_lane30_strm0_tmp     ;
  reg [31:0] pe9_lane30_strm1 [0:4095];
  reg [31:0] pe9_lane30_strm1_tmp     ;
  reg [31:0] pe9_lane31_strm0 [0:4095];
  reg [31:0] pe9_lane31_strm0_tmp     ;
  reg [31:0] pe9_lane31_strm1 [0:4095];
  reg [31:0] pe9_lane31_strm1_tmp     ;
  reg [31:0] pe10_lane0_strm0 [0:4095];
  reg [31:0] pe10_lane0_strm0_tmp     ;
  reg [31:0] pe10_lane0_strm1 [0:4095];
  reg [31:0] pe10_lane0_strm1_tmp     ;
  reg [31:0] pe10_lane1_strm0 [0:4095];
  reg [31:0] pe10_lane1_strm0_tmp     ;
  reg [31:0] pe10_lane1_strm1 [0:4095];
  reg [31:0] pe10_lane1_strm1_tmp     ;
  reg [31:0] pe10_lane2_strm0 [0:4095];
  reg [31:0] pe10_lane2_strm0_tmp     ;
  reg [31:0] pe10_lane2_strm1 [0:4095];
  reg [31:0] pe10_lane2_strm1_tmp     ;
  reg [31:0] pe10_lane3_strm0 [0:4095];
  reg [31:0] pe10_lane3_strm0_tmp     ;
  reg [31:0] pe10_lane3_strm1 [0:4095];
  reg [31:0] pe10_lane3_strm1_tmp     ;
  reg [31:0] pe10_lane4_strm0 [0:4095];
  reg [31:0] pe10_lane4_strm0_tmp     ;
  reg [31:0] pe10_lane4_strm1 [0:4095];
  reg [31:0] pe10_lane4_strm1_tmp     ;
  reg [31:0] pe10_lane5_strm0 [0:4095];
  reg [31:0] pe10_lane5_strm0_tmp     ;
  reg [31:0] pe10_lane5_strm1 [0:4095];
  reg [31:0] pe10_lane5_strm1_tmp     ;
  reg [31:0] pe10_lane6_strm0 [0:4095];
  reg [31:0] pe10_lane6_strm0_tmp     ;
  reg [31:0] pe10_lane6_strm1 [0:4095];
  reg [31:0] pe10_lane6_strm1_tmp     ;
  reg [31:0] pe10_lane7_strm0 [0:4095];
  reg [31:0] pe10_lane7_strm0_tmp     ;
  reg [31:0] pe10_lane7_strm1 [0:4095];
  reg [31:0] pe10_lane7_strm1_tmp     ;
  reg [31:0] pe10_lane8_strm0 [0:4095];
  reg [31:0] pe10_lane8_strm0_tmp     ;
  reg [31:0] pe10_lane8_strm1 [0:4095];
  reg [31:0] pe10_lane8_strm1_tmp     ;
  reg [31:0] pe10_lane9_strm0 [0:4095];
  reg [31:0] pe10_lane9_strm0_tmp     ;
  reg [31:0] pe10_lane9_strm1 [0:4095];
  reg [31:0] pe10_lane9_strm1_tmp     ;
  reg [31:0] pe10_lane10_strm0 [0:4095];
  reg [31:0] pe10_lane10_strm0_tmp     ;
  reg [31:0] pe10_lane10_strm1 [0:4095];
  reg [31:0] pe10_lane10_strm1_tmp     ;
  reg [31:0] pe10_lane11_strm0 [0:4095];
  reg [31:0] pe10_lane11_strm0_tmp     ;
  reg [31:0] pe10_lane11_strm1 [0:4095];
  reg [31:0] pe10_lane11_strm1_tmp     ;
  reg [31:0] pe10_lane12_strm0 [0:4095];
  reg [31:0] pe10_lane12_strm0_tmp     ;
  reg [31:0] pe10_lane12_strm1 [0:4095];
  reg [31:0] pe10_lane12_strm1_tmp     ;
  reg [31:0] pe10_lane13_strm0 [0:4095];
  reg [31:0] pe10_lane13_strm0_tmp     ;
  reg [31:0] pe10_lane13_strm1 [0:4095];
  reg [31:0] pe10_lane13_strm1_tmp     ;
  reg [31:0] pe10_lane14_strm0 [0:4095];
  reg [31:0] pe10_lane14_strm0_tmp     ;
  reg [31:0] pe10_lane14_strm1 [0:4095];
  reg [31:0] pe10_lane14_strm1_tmp     ;
  reg [31:0] pe10_lane15_strm0 [0:4095];
  reg [31:0] pe10_lane15_strm0_tmp     ;
  reg [31:0] pe10_lane15_strm1 [0:4095];
  reg [31:0] pe10_lane15_strm1_tmp     ;
  reg [31:0] pe10_lane16_strm0 [0:4095];
  reg [31:0] pe10_lane16_strm0_tmp     ;
  reg [31:0] pe10_lane16_strm1 [0:4095];
  reg [31:0] pe10_lane16_strm1_tmp     ;
  reg [31:0] pe10_lane17_strm0 [0:4095];
  reg [31:0] pe10_lane17_strm0_tmp     ;
  reg [31:0] pe10_lane17_strm1 [0:4095];
  reg [31:0] pe10_lane17_strm1_tmp     ;
  reg [31:0] pe10_lane18_strm0 [0:4095];
  reg [31:0] pe10_lane18_strm0_tmp     ;
  reg [31:0] pe10_lane18_strm1 [0:4095];
  reg [31:0] pe10_lane18_strm1_tmp     ;
  reg [31:0] pe10_lane19_strm0 [0:4095];
  reg [31:0] pe10_lane19_strm0_tmp     ;
  reg [31:0] pe10_lane19_strm1 [0:4095];
  reg [31:0] pe10_lane19_strm1_tmp     ;
  reg [31:0] pe10_lane20_strm0 [0:4095];
  reg [31:0] pe10_lane20_strm0_tmp     ;
  reg [31:0] pe10_lane20_strm1 [0:4095];
  reg [31:0] pe10_lane20_strm1_tmp     ;
  reg [31:0] pe10_lane21_strm0 [0:4095];
  reg [31:0] pe10_lane21_strm0_tmp     ;
  reg [31:0] pe10_lane21_strm1 [0:4095];
  reg [31:0] pe10_lane21_strm1_tmp     ;
  reg [31:0] pe10_lane22_strm0 [0:4095];
  reg [31:0] pe10_lane22_strm0_tmp     ;
  reg [31:0] pe10_lane22_strm1 [0:4095];
  reg [31:0] pe10_lane22_strm1_tmp     ;
  reg [31:0] pe10_lane23_strm0 [0:4095];
  reg [31:0] pe10_lane23_strm0_tmp     ;
  reg [31:0] pe10_lane23_strm1 [0:4095];
  reg [31:0] pe10_lane23_strm1_tmp     ;
  reg [31:0] pe10_lane24_strm0 [0:4095];
  reg [31:0] pe10_lane24_strm0_tmp     ;
  reg [31:0] pe10_lane24_strm1 [0:4095];
  reg [31:0] pe10_lane24_strm1_tmp     ;
  reg [31:0] pe10_lane25_strm0 [0:4095];
  reg [31:0] pe10_lane25_strm0_tmp     ;
  reg [31:0] pe10_lane25_strm1 [0:4095];
  reg [31:0] pe10_lane25_strm1_tmp     ;
  reg [31:0] pe10_lane26_strm0 [0:4095];
  reg [31:0] pe10_lane26_strm0_tmp     ;
  reg [31:0] pe10_lane26_strm1 [0:4095];
  reg [31:0] pe10_lane26_strm1_tmp     ;
  reg [31:0] pe10_lane27_strm0 [0:4095];
  reg [31:0] pe10_lane27_strm0_tmp     ;
  reg [31:0] pe10_lane27_strm1 [0:4095];
  reg [31:0] pe10_lane27_strm1_tmp     ;
  reg [31:0] pe10_lane28_strm0 [0:4095];
  reg [31:0] pe10_lane28_strm0_tmp     ;
  reg [31:0] pe10_lane28_strm1 [0:4095];
  reg [31:0] pe10_lane28_strm1_tmp     ;
  reg [31:0] pe10_lane29_strm0 [0:4095];
  reg [31:0] pe10_lane29_strm0_tmp     ;
  reg [31:0] pe10_lane29_strm1 [0:4095];
  reg [31:0] pe10_lane29_strm1_tmp     ;
  reg [31:0] pe10_lane30_strm0 [0:4095];
  reg [31:0] pe10_lane30_strm0_tmp     ;
  reg [31:0] pe10_lane30_strm1 [0:4095];
  reg [31:0] pe10_lane30_strm1_tmp     ;
  reg [31:0] pe10_lane31_strm0 [0:4095];
  reg [31:0] pe10_lane31_strm0_tmp     ;
  reg [31:0] pe10_lane31_strm1 [0:4095];
  reg [31:0] pe10_lane31_strm1_tmp     ;
  reg [31:0] pe11_lane0_strm0 [0:4095];
  reg [31:0] pe11_lane0_strm0_tmp     ;
  reg [31:0] pe11_lane0_strm1 [0:4095];
  reg [31:0] pe11_lane0_strm1_tmp     ;
  reg [31:0] pe11_lane1_strm0 [0:4095];
  reg [31:0] pe11_lane1_strm0_tmp     ;
  reg [31:0] pe11_lane1_strm1 [0:4095];
  reg [31:0] pe11_lane1_strm1_tmp     ;
  reg [31:0] pe11_lane2_strm0 [0:4095];
  reg [31:0] pe11_lane2_strm0_tmp     ;
  reg [31:0] pe11_lane2_strm1 [0:4095];
  reg [31:0] pe11_lane2_strm1_tmp     ;
  reg [31:0] pe11_lane3_strm0 [0:4095];
  reg [31:0] pe11_lane3_strm0_tmp     ;
  reg [31:0] pe11_lane3_strm1 [0:4095];
  reg [31:0] pe11_lane3_strm1_tmp     ;
  reg [31:0] pe11_lane4_strm0 [0:4095];
  reg [31:0] pe11_lane4_strm0_tmp     ;
  reg [31:0] pe11_lane4_strm1 [0:4095];
  reg [31:0] pe11_lane4_strm1_tmp     ;
  reg [31:0] pe11_lane5_strm0 [0:4095];
  reg [31:0] pe11_lane5_strm0_tmp     ;
  reg [31:0] pe11_lane5_strm1 [0:4095];
  reg [31:0] pe11_lane5_strm1_tmp     ;
  reg [31:0] pe11_lane6_strm0 [0:4095];
  reg [31:0] pe11_lane6_strm0_tmp     ;
  reg [31:0] pe11_lane6_strm1 [0:4095];
  reg [31:0] pe11_lane6_strm1_tmp     ;
  reg [31:0] pe11_lane7_strm0 [0:4095];
  reg [31:0] pe11_lane7_strm0_tmp     ;
  reg [31:0] pe11_lane7_strm1 [0:4095];
  reg [31:0] pe11_lane7_strm1_tmp     ;
  reg [31:0] pe11_lane8_strm0 [0:4095];
  reg [31:0] pe11_lane8_strm0_tmp     ;
  reg [31:0] pe11_lane8_strm1 [0:4095];
  reg [31:0] pe11_lane8_strm1_tmp     ;
  reg [31:0] pe11_lane9_strm0 [0:4095];
  reg [31:0] pe11_lane9_strm0_tmp     ;
  reg [31:0] pe11_lane9_strm1 [0:4095];
  reg [31:0] pe11_lane9_strm1_tmp     ;
  reg [31:0] pe11_lane10_strm0 [0:4095];
  reg [31:0] pe11_lane10_strm0_tmp     ;
  reg [31:0] pe11_lane10_strm1 [0:4095];
  reg [31:0] pe11_lane10_strm1_tmp     ;
  reg [31:0] pe11_lane11_strm0 [0:4095];
  reg [31:0] pe11_lane11_strm0_tmp     ;
  reg [31:0] pe11_lane11_strm1 [0:4095];
  reg [31:0] pe11_lane11_strm1_tmp     ;
  reg [31:0] pe11_lane12_strm0 [0:4095];
  reg [31:0] pe11_lane12_strm0_tmp     ;
  reg [31:0] pe11_lane12_strm1 [0:4095];
  reg [31:0] pe11_lane12_strm1_tmp     ;
  reg [31:0] pe11_lane13_strm0 [0:4095];
  reg [31:0] pe11_lane13_strm0_tmp     ;
  reg [31:0] pe11_lane13_strm1 [0:4095];
  reg [31:0] pe11_lane13_strm1_tmp     ;
  reg [31:0] pe11_lane14_strm0 [0:4095];
  reg [31:0] pe11_lane14_strm0_tmp     ;
  reg [31:0] pe11_lane14_strm1 [0:4095];
  reg [31:0] pe11_lane14_strm1_tmp     ;
  reg [31:0] pe11_lane15_strm0 [0:4095];
  reg [31:0] pe11_lane15_strm0_tmp     ;
  reg [31:0] pe11_lane15_strm1 [0:4095];
  reg [31:0] pe11_lane15_strm1_tmp     ;
  reg [31:0] pe11_lane16_strm0 [0:4095];
  reg [31:0] pe11_lane16_strm0_tmp     ;
  reg [31:0] pe11_lane16_strm1 [0:4095];
  reg [31:0] pe11_lane16_strm1_tmp     ;
  reg [31:0] pe11_lane17_strm0 [0:4095];
  reg [31:0] pe11_lane17_strm0_tmp     ;
  reg [31:0] pe11_lane17_strm1 [0:4095];
  reg [31:0] pe11_lane17_strm1_tmp     ;
  reg [31:0] pe11_lane18_strm0 [0:4095];
  reg [31:0] pe11_lane18_strm0_tmp     ;
  reg [31:0] pe11_lane18_strm1 [0:4095];
  reg [31:0] pe11_lane18_strm1_tmp     ;
  reg [31:0] pe11_lane19_strm0 [0:4095];
  reg [31:0] pe11_lane19_strm0_tmp     ;
  reg [31:0] pe11_lane19_strm1 [0:4095];
  reg [31:0] pe11_lane19_strm1_tmp     ;
  reg [31:0] pe11_lane20_strm0 [0:4095];
  reg [31:0] pe11_lane20_strm0_tmp     ;
  reg [31:0] pe11_lane20_strm1 [0:4095];
  reg [31:0] pe11_lane20_strm1_tmp     ;
  reg [31:0] pe11_lane21_strm0 [0:4095];
  reg [31:0] pe11_lane21_strm0_tmp     ;
  reg [31:0] pe11_lane21_strm1 [0:4095];
  reg [31:0] pe11_lane21_strm1_tmp     ;
  reg [31:0] pe11_lane22_strm0 [0:4095];
  reg [31:0] pe11_lane22_strm0_tmp     ;
  reg [31:0] pe11_lane22_strm1 [0:4095];
  reg [31:0] pe11_lane22_strm1_tmp     ;
  reg [31:0] pe11_lane23_strm0 [0:4095];
  reg [31:0] pe11_lane23_strm0_tmp     ;
  reg [31:0] pe11_lane23_strm1 [0:4095];
  reg [31:0] pe11_lane23_strm1_tmp     ;
  reg [31:0] pe11_lane24_strm0 [0:4095];
  reg [31:0] pe11_lane24_strm0_tmp     ;
  reg [31:0] pe11_lane24_strm1 [0:4095];
  reg [31:0] pe11_lane24_strm1_tmp     ;
  reg [31:0] pe11_lane25_strm0 [0:4095];
  reg [31:0] pe11_lane25_strm0_tmp     ;
  reg [31:0] pe11_lane25_strm1 [0:4095];
  reg [31:0] pe11_lane25_strm1_tmp     ;
  reg [31:0] pe11_lane26_strm0 [0:4095];
  reg [31:0] pe11_lane26_strm0_tmp     ;
  reg [31:0] pe11_lane26_strm1 [0:4095];
  reg [31:0] pe11_lane26_strm1_tmp     ;
  reg [31:0] pe11_lane27_strm0 [0:4095];
  reg [31:0] pe11_lane27_strm0_tmp     ;
  reg [31:0] pe11_lane27_strm1 [0:4095];
  reg [31:0] pe11_lane27_strm1_tmp     ;
  reg [31:0] pe11_lane28_strm0 [0:4095];
  reg [31:0] pe11_lane28_strm0_tmp     ;
  reg [31:0] pe11_lane28_strm1 [0:4095];
  reg [31:0] pe11_lane28_strm1_tmp     ;
  reg [31:0] pe11_lane29_strm0 [0:4095];
  reg [31:0] pe11_lane29_strm0_tmp     ;
  reg [31:0] pe11_lane29_strm1 [0:4095];
  reg [31:0] pe11_lane29_strm1_tmp     ;
  reg [31:0] pe11_lane30_strm0 [0:4095];
  reg [31:0] pe11_lane30_strm0_tmp     ;
  reg [31:0] pe11_lane30_strm1 [0:4095];
  reg [31:0] pe11_lane30_strm1_tmp     ;
  reg [31:0] pe11_lane31_strm0 [0:4095];
  reg [31:0] pe11_lane31_strm0_tmp     ;
  reg [31:0] pe11_lane31_strm1 [0:4095];
  reg [31:0] pe11_lane31_strm1_tmp     ;
  reg [31:0] pe12_lane0_strm0 [0:4095];
  reg [31:0] pe12_lane0_strm0_tmp     ;
  reg [31:0] pe12_lane0_strm1 [0:4095];
  reg [31:0] pe12_lane0_strm1_tmp     ;
  reg [31:0] pe12_lane1_strm0 [0:4095];
  reg [31:0] pe12_lane1_strm0_tmp     ;
  reg [31:0] pe12_lane1_strm1 [0:4095];
  reg [31:0] pe12_lane1_strm1_tmp     ;
  reg [31:0] pe12_lane2_strm0 [0:4095];
  reg [31:0] pe12_lane2_strm0_tmp     ;
  reg [31:0] pe12_lane2_strm1 [0:4095];
  reg [31:0] pe12_lane2_strm1_tmp     ;
  reg [31:0] pe12_lane3_strm0 [0:4095];
  reg [31:0] pe12_lane3_strm0_tmp     ;
  reg [31:0] pe12_lane3_strm1 [0:4095];
  reg [31:0] pe12_lane3_strm1_tmp     ;
  reg [31:0] pe12_lane4_strm0 [0:4095];
  reg [31:0] pe12_lane4_strm0_tmp     ;
  reg [31:0] pe12_lane4_strm1 [0:4095];
  reg [31:0] pe12_lane4_strm1_tmp     ;
  reg [31:0] pe12_lane5_strm0 [0:4095];
  reg [31:0] pe12_lane5_strm0_tmp     ;
  reg [31:0] pe12_lane5_strm1 [0:4095];
  reg [31:0] pe12_lane5_strm1_tmp     ;
  reg [31:0] pe12_lane6_strm0 [0:4095];
  reg [31:0] pe12_lane6_strm0_tmp     ;
  reg [31:0] pe12_lane6_strm1 [0:4095];
  reg [31:0] pe12_lane6_strm1_tmp     ;
  reg [31:0] pe12_lane7_strm0 [0:4095];
  reg [31:0] pe12_lane7_strm0_tmp     ;
  reg [31:0] pe12_lane7_strm1 [0:4095];
  reg [31:0] pe12_lane7_strm1_tmp     ;
  reg [31:0] pe12_lane8_strm0 [0:4095];
  reg [31:0] pe12_lane8_strm0_tmp     ;
  reg [31:0] pe12_lane8_strm1 [0:4095];
  reg [31:0] pe12_lane8_strm1_tmp     ;
  reg [31:0] pe12_lane9_strm0 [0:4095];
  reg [31:0] pe12_lane9_strm0_tmp     ;
  reg [31:0] pe12_lane9_strm1 [0:4095];
  reg [31:0] pe12_lane9_strm1_tmp     ;
  reg [31:0] pe12_lane10_strm0 [0:4095];
  reg [31:0] pe12_lane10_strm0_tmp     ;
  reg [31:0] pe12_lane10_strm1 [0:4095];
  reg [31:0] pe12_lane10_strm1_tmp     ;
  reg [31:0] pe12_lane11_strm0 [0:4095];
  reg [31:0] pe12_lane11_strm0_tmp     ;
  reg [31:0] pe12_lane11_strm1 [0:4095];
  reg [31:0] pe12_lane11_strm1_tmp     ;
  reg [31:0] pe12_lane12_strm0 [0:4095];
  reg [31:0] pe12_lane12_strm0_tmp     ;
  reg [31:0] pe12_lane12_strm1 [0:4095];
  reg [31:0] pe12_lane12_strm1_tmp     ;
  reg [31:0] pe12_lane13_strm0 [0:4095];
  reg [31:0] pe12_lane13_strm0_tmp     ;
  reg [31:0] pe12_lane13_strm1 [0:4095];
  reg [31:0] pe12_lane13_strm1_tmp     ;
  reg [31:0] pe12_lane14_strm0 [0:4095];
  reg [31:0] pe12_lane14_strm0_tmp     ;
  reg [31:0] pe12_lane14_strm1 [0:4095];
  reg [31:0] pe12_lane14_strm1_tmp     ;
  reg [31:0] pe12_lane15_strm0 [0:4095];
  reg [31:0] pe12_lane15_strm0_tmp     ;
  reg [31:0] pe12_lane15_strm1 [0:4095];
  reg [31:0] pe12_lane15_strm1_tmp     ;
  reg [31:0] pe12_lane16_strm0 [0:4095];
  reg [31:0] pe12_lane16_strm0_tmp     ;
  reg [31:0] pe12_lane16_strm1 [0:4095];
  reg [31:0] pe12_lane16_strm1_tmp     ;
  reg [31:0] pe12_lane17_strm0 [0:4095];
  reg [31:0] pe12_lane17_strm0_tmp     ;
  reg [31:0] pe12_lane17_strm1 [0:4095];
  reg [31:0] pe12_lane17_strm1_tmp     ;
  reg [31:0] pe12_lane18_strm0 [0:4095];
  reg [31:0] pe12_lane18_strm0_tmp     ;
  reg [31:0] pe12_lane18_strm1 [0:4095];
  reg [31:0] pe12_lane18_strm1_tmp     ;
  reg [31:0] pe12_lane19_strm0 [0:4095];
  reg [31:0] pe12_lane19_strm0_tmp     ;
  reg [31:0] pe12_lane19_strm1 [0:4095];
  reg [31:0] pe12_lane19_strm1_tmp     ;
  reg [31:0] pe12_lane20_strm0 [0:4095];
  reg [31:0] pe12_lane20_strm0_tmp     ;
  reg [31:0] pe12_lane20_strm1 [0:4095];
  reg [31:0] pe12_lane20_strm1_tmp     ;
  reg [31:0] pe12_lane21_strm0 [0:4095];
  reg [31:0] pe12_lane21_strm0_tmp     ;
  reg [31:0] pe12_lane21_strm1 [0:4095];
  reg [31:0] pe12_lane21_strm1_tmp     ;
  reg [31:0] pe12_lane22_strm0 [0:4095];
  reg [31:0] pe12_lane22_strm0_tmp     ;
  reg [31:0] pe12_lane22_strm1 [0:4095];
  reg [31:0] pe12_lane22_strm1_tmp     ;
  reg [31:0] pe12_lane23_strm0 [0:4095];
  reg [31:0] pe12_lane23_strm0_tmp     ;
  reg [31:0] pe12_lane23_strm1 [0:4095];
  reg [31:0] pe12_lane23_strm1_tmp     ;
  reg [31:0] pe12_lane24_strm0 [0:4095];
  reg [31:0] pe12_lane24_strm0_tmp     ;
  reg [31:0] pe12_lane24_strm1 [0:4095];
  reg [31:0] pe12_lane24_strm1_tmp     ;
  reg [31:0] pe12_lane25_strm0 [0:4095];
  reg [31:0] pe12_lane25_strm0_tmp     ;
  reg [31:0] pe12_lane25_strm1 [0:4095];
  reg [31:0] pe12_lane25_strm1_tmp     ;
  reg [31:0] pe12_lane26_strm0 [0:4095];
  reg [31:0] pe12_lane26_strm0_tmp     ;
  reg [31:0] pe12_lane26_strm1 [0:4095];
  reg [31:0] pe12_lane26_strm1_tmp     ;
  reg [31:0] pe12_lane27_strm0 [0:4095];
  reg [31:0] pe12_lane27_strm0_tmp     ;
  reg [31:0] pe12_lane27_strm1 [0:4095];
  reg [31:0] pe12_lane27_strm1_tmp     ;
  reg [31:0] pe12_lane28_strm0 [0:4095];
  reg [31:0] pe12_lane28_strm0_tmp     ;
  reg [31:0] pe12_lane28_strm1 [0:4095];
  reg [31:0] pe12_lane28_strm1_tmp     ;
  reg [31:0] pe12_lane29_strm0 [0:4095];
  reg [31:0] pe12_lane29_strm0_tmp     ;
  reg [31:0] pe12_lane29_strm1 [0:4095];
  reg [31:0] pe12_lane29_strm1_tmp     ;
  reg [31:0] pe12_lane30_strm0 [0:4095];
  reg [31:0] pe12_lane30_strm0_tmp     ;
  reg [31:0] pe12_lane30_strm1 [0:4095];
  reg [31:0] pe12_lane30_strm1_tmp     ;
  reg [31:0] pe12_lane31_strm0 [0:4095];
  reg [31:0] pe12_lane31_strm0_tmp     ;
  reg [31:0] pe12_lane31_strm1 [0:4095];
  reg [31:0] pe12_lane31_strm1_tmp     ;
  reg [31:0] pe13_lane0_strm0 [0:4095];
  reg [31:0] pe13_lane0_strm0_tmp     ;
  reg [31:0] pe13_lane0_strm1 [0:4095];
  reg [31:0] pe13_lane0_strm1_tmp     ;
  reg [31:0] pe13_lane1_strm0 [0:4095];
  reg [31:0] pe13_lane1_strm0_tmp     ;
  reg [31:0] pe13_lane1_strm1 [0:4095];
  reg [31:0] pe13_lane1_strm1_tmp     ;
  reg [31:0] pe13_lane2_strm0 [0:4095];
  reg [31:0] pe13_lane2_strm0_tmp     ;
  reg [31:0] pe13_lane2_strm1 [0:4095];
  reg [31:0] pe13_lane2_strm1_tmp     ;
  reg [31:0] pe13_lane3_strm0 [0:4095];
  reg [31:0] pe13_lane3_strm0_tmp     ;
  reg [31:0] pe13_lane3_strm1 [0:4095];
  reg [31:0] pe13_lane3_strm1_tmp     ;
  reg [31:0] pe13_lane4_strm0 [0:4095];
  reg [31:0] pe13_lane4_strm0_tmp     ;
  reg [31:0] pe13_lane4_strm1 [0:4095];
  reg [31:0] pe13_lane4_strm1_tmp     ;
  reg [31:0] pe13_lane5_strm0 [0:4095];
  reg [31:0] pe13_lane5_strm0_tmp     ;
  reg [31:0] pe13_lane5_strm1 [0:4095];
  reg [31:0] pe13_lane5_strm1_tmp     ;
  reg [31:0] pe13_lane6_strm0 [0:4095];
  reg [31:0] pe13_lane6_strm0_tmp     ;
  reg [31:0] pe13_lane6_strm1 [0:4095];
  reg [31:0] pe13_lane6_strm1_tmp     ;
  reg [31:0] pe13_lane7_strm0 [0:4095];
  reg [31:0] pe13_lane7_strm0_tmp     ;
  reg [31:0] pe13_lane7_strm1 [0:4095];
  reg [31:0] pe13_lane7_strm1_tmp     ;
  reg [31:0] pe13_lane8_strm0 [0:4095];
  reg [31:0] pe13_lane8_strm0_tmp     ;
  reg [31:0] pe13_lane8_strm1 [0:4095];
  reg [31:0] pe13_lane8_strm1_tmp     ;
  reg [31:0] pe13_lane9_strm0 [0:4095];
  reg [31:0] pe13_lane9_strm0_tmp     ;
  reg [31:0] pe13_lane9_strm1 [0:4095];
  reg [31:0] pe13_lane9_strm1_tmp     ;
  reg [31:0] pe13_lane10_strm0 [0:4095];
  reg [31:0] pe13_lane10_strm0_tmp     ;
  reg [31:0] pe13_lane10_strm1 [0:4095];
  reg [31:0] pe13_lane10_strm1_tmp     ;
  reg [31:0] pe13_lane11_strm0 [0:4095];
  reg [31:0] pe13_lane11_strm0_tmp     ;
  reg [31:0] pe13_lane11_strm1 [0:4095];
  reg [31:0] pe13_lane11_strm1_tmp     ;
  reg [31:0] pe13_lane12_strm0 [0:4095];
  reg [31:0] pe13_lane12_strm0_tmp     ;
  reg [31:0] pe13_lane12_strm1 [0:4095];
  reg [31:0] pe13_lane12_strm1_tmp     ;
  reg [31:0] pe13_lane13_strm0 [0:4095];
  reg [31:0] pe13_lane13_strm0_tmp     ;
  reg [31:0] pe13_lane13_strm1 [0:4095];
  reg [31:0] pe13_lane13_strm1_tmp     ;
  reg [31:0] pe13_lane14_strm0 [0:4095];
  reg [31:0] pe13_lane14_strm0_tmp     ;
  reg [31:0] pe13_lane14_strm1 [0:4095];
  reg [31:0] pe13_lane14_strm1_tmp     ;
  reg [31:0] pe13_lane15_strm0 [0:4095];
  reg [31:0] pe13_lane15_strm0_tmp     ;
  reg [31:0] pe13_lane15_strm1 [0:4095];
  reg [31:0] pe13_lane15_strm1_tmp     ;
  reg [31:0] pe13_lane16_strm0 [0:4095];
  reg [31:0] pe13_lane16_strm0_tmp     ;
  reg [31:0] pe13_lane16_strm1 [0:4095];
  reg [31:0] pe13_lane16_strm1_tmp     ;
  reg [31:0] pe13_lane17_strm0 [0:4095];
  reg [31:0] pe13_lane17_strm0_tmp     ;
  reg [31:0] pe13_lane17_strm1 [0:4095];
  reg [31:0] pe13_lane17_strm1_tmp     ;
  reg [31:0] pe13_lane18_strm0 [0:4095];
  reg [31:0] pe13_lane18_strm0_tmp     ;
  reg [31:0] pe13_lane18_strm1 [0:4095];
  reg [31:0] pe13_lane18_strm1_tmp     ;
  reg [31:0] pe13_lane19_strm0 [0:4095];
  reg [31:0] pe13_lane19_strm0_tmp     ;
  reg [31:0] pe13_lane19_strm1 [0:4095];
  reg [31:0] pe13_lane19_strm1_tmp     ;
  reg [31:0] pe13_lane20_strm0 [0:4095];
  reg [31:0] pe13_lane20_strm0_tmp     ;
  reg [31:0] pe13_lane20_strm1 [0:4095];
  reg [31:0] pe13_lane20_strm1_tmp     ;
  reg [31:0] pe13_lane21_strm0 [0:4095];
  reg [31:0] pe13_lane21_strm0_tmp     ;
  reg [31:0] pe13_lane21_strm1 [0:4095];
  reg [31:0] pe13_lane21_strm1_tmp     ;
  reg [31:0] pe13_lane22_strm0 [0:4095];
  reg [31:0] pe13_lane22_strm0_tmp     ;
  reg [31:0] pe13_lane22_strm1 [0:4095];
  reg [31:0] pe13_lane22_strm1_tmp     ;
  reg [31:0] pe13_lane23_strm0 [0:4095];
  reg [31:0] pe13_lane23_strm0_tmp     ;
  reg [31:0] pe13_lane23_strm1 [0:4095];
  reg [31:0] pe13_lane23_strm1_tmp     ;
  reg [31:0] pe13_lane24_strm0 [0:4095];
  reg [31:0] pe13_lane24_strm0_tmp     ;
  reg [31:0] pe13_lane24_strm1 [0:4095];
  reg [31:0] pe13_lane24_strm1_tmp     ;
  reg [31:0] pe13_lane25_strm0 [0:4095];
  reg [31:0] pe13_lane25_strm0_tmp     ;
  reg [31:0] pe13_lane25_strm1 [0:4095];
  reg [31:0] pe13_lane25_strm1_tmp     ;
  reg [31:0] pe13_lane26_strm0 [0:4095];
  reg [31:0] pe13_lane26_strm0_tmp     ;
  reg [31:0] pe13_lane26_strm1 [0:4095];
  reg [31:0] pe13_lane26_strm1_tmp     ;
  reg [31:0] pe13_lane27_strm0 [0:4095];
  reg [31:0] pe13_lane27_strm0_tmp     ;
  reg [31:0] pe13_lane27_strm1 [0:4095];
  reg [31:0] pe13_lane27_strm1_tmp     ;
  reg [31:0] pe13_lane28_strm0 [0:4095];
  reg [31:0] pe13_lane28_strm0_tmp     ;
  reg [31:0] pe13_lane28_strm1 [0:4095];
  reg [31:0] pe13_lane28_strm1_tmp     ;
  reg [31:0] pe13_lane29_strm0 [0:4095];
  reg [31:0] pe13_lane29_strm0_tmp     ;
  reg [31:0] pe13_lane29_strm1 [0:4095];
  reg [31:0] pe13_lane29_strm1_tmp     ;
  reg [31:0] pe13_lane30_strm0 [0:4095];
  reg [31:0] pe13_lane30_strm0_tmp     ;
  reg [31:0] pe13_lane30_strm1 [0:4095];
  reg [31:0] pe13_lane30_strm1_tmp     ;
  reg [31:0] pe13_lane31_strm0 [0:4095];
  reg [31:0] pe13_lane31_strm0_tmp     ;
  reg [31:0] pe13_lane31_strm1 [0:4095];
  reg [31:0] pe13_lane31_strm1_tmp     ;
  reg [31:0] pe14_lane0_strm0 [0:4095];
  reg [31:0] pe14_lane0_strm0_tmp     ;
  reg [31:0] pe14_lane0_strm1 [0:4095];
  reg [31:0] pe14_lane0_strm1_tmp     ;
  reg [31:0] pe14_lane1_strm0 [0:4095];
  reg [31:0] pe14_lane1_strm0_tmp     ;
  reg [31:0] pe14_lane1_strm1 [0:4095];
  reg [31:0] pe14_lane1_strm1_tmp     ;
  reg [31:0] pe14_lane2_strm0 [0:4095];
  reg [31:0] pe14_lane2_strm0_tmp     ;
  reg [31:0] pe14_lane2_strm1 [0:4095];
  reg [31:0] pe14_lane2_strm1_tmp     ;
  reg [31:0] pe14_lane3_strm0 [0:4095];
  reg [31:0] pe14_lane3_strm0_tmp     ;
  reg [31:0] pe14_lane3_strm1 [0:4095];
  reg [31:0] pe14_lane3_strm1_tmp     ;
  reg [31:0] pe14_lane4_strm0 [0:4095];
  reg [31:0] pe14_lane4_strm0_tmp     ;
  reg [31:0] pe14_lane4_strm1 [0:4095];
  reg [31:0] pe14_lane4_strm1_tmp     ;
  reg [31:0] pe14_lane5_strm0 [0:4095];
  reg [31:0] pe14_lane5_strm0_tmp     ;
  reg [31:0] pe14_lane5_strm1 [0:4095];
  reg [31:0] pe14_lane5_strm1_tmp     ;
  reg [31:0] pe14_lane6_strm0 [0:4095];
  reg [31:0] pe14_lane6_strm0_tmp     ;
  reg [31:0] pe14_lane6_strm1 [0:4095];
  reg [31:0] pe14_lane6_strm1_tmp     ;
  reg [31:0] pe14_lane7_strm0 [0:4095];
  reg [31:0] pe14_lane7_strm0_tmp     ;
  reg [31:0] pe14_lane7_strm1 [0:4095];
  reg [31:0] pe14_lane7_strm1_tmp     ;
  reg [31:0] pe14_lane8_strm0 [0:4095];
  reg [31:0] pe14_lane8_strm0_tmp     ;
  reg [31:0] pe14_lane8_strm1 [0:4095];
  reg [31:0] pe14_lane8_strm1_tmp     ;
  reg [31:0] pe14_lane9_strm0 [0:4095];
  reg [31:0] pe14_lane9_strm0_tmp     ;
  reg [31:0] pe14_lane9_strm1 [0:4095];
  reg [31:0] pe14_lane9_strm1_tmp     ;
  reg [31:0] pe14_lane10_strm0 [0:4095];
  reg [31:0] pe14_lane10_strm0_tmp     ;
  reg [31:0] pe14_lane10_strm1 [0:4095];
  reg [31:0] pe14_lane10_strm1_tmp     ;
  reg [31:0] pe14_lane11_strm0 [0:4095];
  reg [31:0] pe14_lane11_strm0_tmp     ;
  reg [31:0] pe14_lane11_strm1 [0:4095];
  reg [31:0] pe14_lane11_strm1_tmp     ;
  reg [31:0] pe14_lane12_strm0 [0:4095];
  reg [31:0] pe14_lane12_strm0_tmp     ;
  reg [31:0] pe14_lane12_strm1 [0:4095];
  reg [31:0] pe14_lane12_strm1_tmp     ;
  reg [31:0] pe14_lane13_strm0 [0:4095];
  reg [31:0] pe14_lane13_strm0_tmp     ;
  reg [31:0] pe14_lane13_strm1 [0:4095];
  reg [31:0] pe14_lane13_strm1_tmp     ;
  reg [31:0] pe14_lane14_strm0 [0:4095];
  reg [31:0] pe14_lane14_strm0_tmp     ;
  reg [31:0] pe14_lane14_strm1 [0:4095];
  reg [31:0] pe14_lane14_strm1_tmp     ;
  reg [31:0] pe14_lane15_strm0 [0:4095];
  reg [31:0] pe14_lane15_strm0_tmp     ;
  reg [31:0] pe14_lane15_strm1 [0:4095];
  reg [31:0] pe14_lane15_strm1_tmp     ;
  reg [31:0] pe14_lane16_strm0 [0:4095];
  reg [31:0] pe14_lane16_strm0_tmp     ;
  reg [31:0] pe14_lane16_strm1 [0:4095];
  reg [31:0] pe14_lane16_strm1_tmp     ;
  reg [31:0] pe14_lane17_strm0 [0:4095];
  reg [31:0] pe14_lane17_strm0_tmp     ;
  reg [31:0] pe14_lane17_strm1 [0:4095];
  reg [31:0] pe14_lane17_strm1_tmp     ;
  reg [31:0] pe14_lane18_strm0 [0:4095];
  reg [31:0] pe14_lane18_strm0_tmp     ;
  reg [31:0] pe14_lane18_strm1 [0:4095];
  reg [31:0] pe14_lane18_strm1_tmp     ;
  reg [31:0] pe14_lane19_strm0 [0:4095];
  reg [31:0] pe14_lane19_strm0_tmp     ;
  reg [31:0] pe14_lane19_strm1 [0:4095];
  reg [31:0] pe14_lane19_strm1_tmp     ;
  reg [31:0] pe14_lane20_strm0 [0:4095];
  reg [31:0] pe14_lane20_strm0_tmp     ;
  reg [31:0] pe14_lane20_strm1 [0:4095];
  reg [31:0] pe14_lane20_strm1_tmp     ;
  reg [31:0] pe14_lane21_strm0 [0:4095];
  reg [31:0] pe14_lane21_strm0_tmp     ;
  reg [31:0] pe14_lane21_strm1 [0:4095];
  reg [31:0] pe14_lane21_strm1_tmp     ;
  reg [31:0] pe14_lane22_strm0 [0:4095];
  reg [31:0] pe14_lane22_strm0_tmp     ;
  reg [31:0] pe14_lane22_strm1 [0:4095];
  reg [31:0] pe14_lane22_strm1_tmp     ;
  reg [31:0] pe14_lane23_strm0 [0:4095];
  reg [31:0] pe14_lane23_strm0_tmp     ;
  reg [31:0] pe14_lane23_strm1 [0:4095];
  reg [31:0] pe14_lane23_strm1_tmp     ;
  reg [31:0] pe14_lane24_strm0 [0:4095];
  reg [31:0] pe14_lane24_strm0_tmp     ;
  reg [31:0] pe14_lane24_strm1 [0:4095];
  reg [31:0] pe14_lane24_strm1_tmp     ;
  reg [31:0] pe14_lane25_strm0 [0:4095];
  reg [31:0] pe14_lane25_strm0_tmp     ;
  reg [31:0] pe14_lane25_strm1 [0:4095];
  reg [31:0] pe14_lane25_strm1_tmp     ;
  reg [31:0] pe14_lane26_strm0 [0:4095];
  reg [31:0] pe14_lane26_strm0_tmp     ;
  reg [31:0] pe14_lane26_strm1 [0:4095];
  reg [31:0] pe14_lane26_strm1_tmp     ;
  reg [31:0] pe14_lane27_strm0 [0:4095];
  reg [31:0] pe14_lane27_strm0_tmp     ;
  reg [31:0] pe14_lane27_strm1 [0:4095];
  reg [31:0] pe14_lane27_strm1_tmp     ;
  reg [31:0] pe14_lane28_strm0 [0:4095];
  reg [31:0] pe14_lane28_strm0_tmp     ;
  reg [31:0] pe14_lane28_strm1 [0:4095];
  reg [31:0] pe14_lane28_strm1_tmp     ;
  reg [31:0] pe14_lane29_strm0 [0:4095];
  reg [31:0] pe14_lane29_strm0_tmp     ;
  reg [31:0] pe14_lane29_strm1 [0:4095];
  reg [31:0] pe14_lane29_strm1_tmp     ;
  reg [31:0] pe14_lane30_strm0 [0:4095];
  reg [31:0] pe14_lane30_strm0_tmp     ;
  reg [31:0] pe14_lane30_strm1 [0:4095];
  reg [31:0] pe14_lane30_strm1_tmp     ;
  reg [31:0] pe14_lane31_strm0 [0:4095];
  reg [31:0] pe14_lane31_strm0_tmp     ;
  reg [31:0] pe14_lane31_strm1 [0:4095];
  reg [31:0] pe14_lane31_strm1_tmp     ;
  reg [31:0] pe15_lane0_strm0 [0:4095];
  reg [31:0] pe15_lane0_strm0_tmp     ;
  reg [31:0] pe15_lane0_strm1 [0:4095];
  reg [31:0] pe15_lane0_strm1_tmp     ;
  reg [31:0] pe15_lane1_strm0 [0:4095];
  reg [31:0] pe15_lane1_strm0_tmp     ;
  reg [31:0] pe15_lane1_strm1 [0:4095];
  reg [31:0] pe15_lane1_strm1_tmp     ;
  reg [31:0] pe15_lane2_strm0 [0:4095];
  reg [31:0] pe15_lane2_strm0_tmp     ;
  reg [31:0] pe15_lane2_strm1 [0:4095];
  reg [31:0] pe15_lane2_strm1_tmp     ;
  reg [31:0] pe15_lane3_strm0 [0:4095];
  reg [31:0] pe15_lane3_strm0_tmp     ;
  reg [31:0] pe15_lane3_strm1 [0:4095];
  reg [31:0] pe15_lane3_strm1_tmp     ;
  reg [31:0] pe15_lane4_strm0 [0:4095];
  reg [31:0] pe15_lane4_strm0_tmp     ;
  reg [31:0] pe15_lane4_strm1 [0:4095];
  reg [31:0] pe15_lane4_strm1_tmp     ;
  reg [31:0] pe15_lane5_strm0 [0:4095];
  reg [31:0] pe15_lane5_strm0_tmp     ;
  reg [31:0] pe15_lane5_strm1 [0:4095];
  reg [31:0] pe15_lane5_strm1_tmp     ;
  reg [31:0] pe15_lane6_strm0 [0:4095];
  reg [31:0] pe15_lane6_strm0_tmp     ;
  reg [31:0] pe15_lane6_strm1 [0:4095];
  reg [31:0] pe15_lane6_strm1_tmp     ;
  reg [31:0] pe15_lane7_strm0 [0:4095];
  reg [31:0] pe15_lane7_strm0_tmp     ;
  reg [31:0] pe15_lane7_strm1 [0:4095];
  reg [31:0] pe15_lane7_strm1_tmp     ;
  reg [31:0] pe15_lane8_strm0 [0:4095];
  reg [31:0] pe15_lane8_strm0_tmp     ;
  reg [31:0] pe15_lane8_strm1 [0:4095];
  reg [31:0] pe15_lane8_strm1_tmp     ;
  reg [31:0] pe15_lane9_strm0 [0:4095];
  reg [31:0] pe15_lane9_strm0_tmp     ;
  reg [31:0] pe15_lane9_strm1 [0:4095];
  reg [31:0] pe15_lane9_strm1_tmp     ;
  reg [31:0] pe15_lane10_strm0 [0:4095];
  reg [31:0] pe15_lane10_strm0_tmp     ;
  reg [31:0] pe15_lane10_strm1 [0:4095];
  reg [31:0] pe15_lane10_strm1_tmp     ;
  reg [31:0] pe15_lane11_strm0 [0:4095];
  reg [31:0] pe15_lane11_strm0_tmp     ;
  reg [31:0] pe15_lane11_strm1 [0:4095];
  reg [31:0] pe15_lane11_strm1_tmp     ;
  reg [31:0] pe15_lane12_strm0 [0:4095];
  reg [31:0] pe15_lane12_strm0_tmp     ;
  reg [31:0] pe15_lane12_strm1 [0:4095];
  reg [31:0] pe15_lane12_strm1_tmp     ;
  reg [31:0] pe15_lane13_strm0 [0:4095];
  reg [31:0] pe15_lane13_strm0_tmp     ;
  reg [31:0] pe15_lane13_strm1 [0:4095];
  reg [31:0] pe15_lane13_strm1_tmp     ;
  reg [31:0] pe15_lane14_strm0 [0:4095];
  reg [31:0] pe15_lane14_strm0_tmp     ;
  reg [31:0] pe15_lane14_strm1 [0:4095];
  reg [31:0] pe15_lane14_strm1_tmp     ;
  reg [31:0] pe15_lane15_strm0 [0:4095];
  reg [31:0] pe15_lane15_strm0_tmp     ;
  reg [31:0] pe15_lane15_strm1 [0:4095];
  reg [31:0] pe15_lane15_strm1_tmp     ;
  reg [31:0] pe15_lane16_strm0 [0:4095];
  reg [31:0] pe15_lane16_strm0_tmp     ;
  reg [31:0] pe15_lane16_strm1 [0:4095];
  reg [31:0] pe15_lane16_strm1_tmp     ;
  reg [31:0] pe15_lane17_strm0 [0:4095];
  reg [31:0] pe15_lane17_strm0_tmp     ;
  reg [31:0] pe15_lane17_strm1 [0:4095];
  reg [31:0] pe15_lane17_strm1_tmp     ;
  reg [31:0] pe15_lane18_strm0 [0:4095];
  reg [31:0] pe15_lane18_strm0_tmp     ;
  reg [31:0] pe15_lane18_strm1 [0:4095];
  reg [31:0] pe15_lane18_strm1_tmp     ;
  reg [31:0] pe15_lane19_strm0 [0:4095];
  reg [31:0] pe15_lane19_strm0_tmp     ;
  reg [31:0] pe15_lane19_strm1 [0:4095];
  reg [31:0] pe15_lane19_strm1_tmp     ;
  reg [31:0] pe15_lane20_strm0 [0:4095];
  reg [31:0] pe15_lane20_strm0_tmp     ;
  reg [31:0] pe15_lane20_strm1 [0:4095];
  reg [31:0] pe15_lane20_strm1_tmp     ;
  reg [31:0] pe15_lane21_strm0 [0:4095];
  reg [31:0] pe15_lane21_strm0_tmp     ;
  reg [31:0] pe15_lane21_strm1 [0:4095];
  reg [31:0] pe15_lane21_strm1_tmp     ;
  reg [31:0] pe15_lane22_strm0 [0:4095];
  reg [31:0] pe15_lane22_strm0_tmp     ;
  reg [31:0] pe15_lane22_strm1 [0:4095];
  reg [31:0] pe15_lane22_strm1_tmp     ;
  reg [31:0] pe15_lane23_strm0 [0:4095];
  reg [31:0] pe15_lane23_strm0_tmp     ;
  reg [31:0] pe15_lane23_strm1 [0:4095];
  reg [31:0] pe15_lane23_strm1_tmp     ;
  reg [31:0] pe15_lane24_strm0 [0:4095];
  reg [31:0] pe15_lane24_strm0_tmp     ;
  reg [31:0] pe15_lane24_strm1 [0:4095];
  reg [31:0] pe15_lane24_strm1_tmp     ;
  reg [31:0] pe15_lane25_strm0 [0:4095];
  reg [31:0] pe15_lane25_strm0_tmp     ;
  reg [31:0] pe15_lane25_strm1 [0:4095];
  reg [31:0] pe15_lane25_strm1_tmp     ;
  reg [31:0] pe15_lane26_strm0 [0:4095];
  reg [31:0] pe15_lane26_strm0_tmp     ;
  reg [31:0] pe15_lane26_strm1 [0:4095];
  reg [31:0] pe15_lane26_strm1_tmp     ;
  reg [31:0] pe15_lane27_strm0 [0:4095];
  reg [31:0] pe15_lane27_strm0_tmp     ;
  reg [31:0] pe15_lane27_strm1 [0:4095];
  reg [31:0] pe15_lane27_strm1_tmp     ;
  reg [31:0] pe15_lane28_strm0 [0:4095];
  reg [31:0] pe15_lane28_strm0_tmp     ;
  reg [31:0] pe15_lane28_strm1 [0:4095];
  reg [31:0] pe15_lane28_strm1_tmp     ;
  reg [31:0] pe15_lane29_strm0 [0:4095];
  reg [31:0] pe15_lane29_strm0_tmp     ;
  reg [31:0] pe15_lane29_strm1 [0:4095];
  reg [31:0] pe15_lane29_strm1_tmp     ;
  reg [31:0] pe15_lane30_strm0 [0:4095];
  reg [31:0] pe15_lane30_strm0_tmp     ;
  reg [31:0] pe15_lane30_strm1 [0:4095];
  reg [31:0] pe15_lane30_strm1_tmp     ;
  reg [31:0] pe15_lane31_strm0 [0:4095];
  reg [31:0] pe15_lane31_strm0_tmp     ;
  reg [31:0] pe15_lane31_strm1 [0:4095];
  reg [31:0] pe15_lane31_strm1_tmp     ;
  reg [31:0] pe16_lane0_strm0 [0:4095];
  reg [31:0] pe16_lane0_strm0_tmp     ;
  reg [31:0] pe16_lane0_strm1 [0:4095];
  reg [31:0] pe16_lane0_strm1_tmp     ;
  reg [31:0] pe16_lane1_strm0 [0:4095];
  reg [31:0] pe16_lane1_strm0_tmp     ;
  reg [31:0] pe16_lane1_strm1 [0:4095];
  reg [31:0] pe16_lane1_strm1_tmp     ;
  reg [31:0] pe16_lane2_strm0 [0:4095];
  reg [31:0] pe16_lane2_strm0_tmp     ;
  reg [31:0] pe16_lane2_strm1 [0:4095];
  reg [31:0] pe16_lane2_strm1_tmp     ;
  reg [31:0] pe16_lane3_strm0 [0:4095];
  reg [31:0] pe16_lane3_strm0_tmp     ;
  reg [31:0] pe16_lane3_strm1 [0:4095];
  reg [31:0] pe16_lane3_strm1_tmp     ;
  reg [31:0] pe16_lane4_strm0 [0:4095];
  reg [31:0] pe16_lane4_strm0_tmp     ;
  reg [31:0] pe16_lane4_strm1 [0:4095];
  reg [31:0] pe16_lane4_strm1_tmp     ;
  reg [31:0] pe16_lane5_strm0 [0:4095];
  reg [31:0] pe16_lane5_strm0_tmp     ;
  reg [31:0] pe16_lane5_strm1 [0:4095];
  reg [31:0] pe16_lane5_strm1_tmp     ;
  reg [31:0] pe16_lane6_strm0 [0:4095];
  reg [31:0] pe16_lane6_strm0_tmp     ;
  reg [31:0] pe16_lane6_strm1 [0:4095];
  reg [31:0] pe16_lane6_strm1_tmp     ;
  reg [31:0] pe16_lane7_strm0 [0:4095];
  reg [31:0] pe16_lane7_strm0_tmp     ;
  reg [31:0] pe16_lane7_strm1 [0:4095];
  reg [31:0] pe16_lane7_strm1_tmp     ;
  reg [31:0] pe16_lane8_strm0 [0:4095];
  reg [31:0] pe16_lane8_strm0_tmp     ;
  reg [31:0] pe16_lane8_strm1 [0:4095];
  reg [31:0] pe16_lane8_strm1_tmp     ;
  reg [31:0] pe16_lane9_strm0 [0:4095];
  reg [31:0] pe16_lane9_strm0_tmp     ;
  reg [31:0] pe16_lane9_strm1 [0:4095];
  reg [31:0] pe16_lane9_strm1_tmp     ;
  reg [31:0] pe16_lane10_strm0 [0:4095];
  reg [31:0] pe16_lane10_strm0_tmp     ;
  reg [31:0] pe16_lane10_strm1 [0:4095];
  reg [31:0] pe16_lane10_strm1_tmp     ;
  reg [31:0] pe16_lane11_strm0 [0:4095];
  reg [31:0] pe16_lane11_strm0_tmp     ;
  reg [31:0] pe16_lane11_strm1 [0:4095];
  reg [31:0] pe16_lane11_strm1_tmp     ;
  reg [31:0] pe16_lane12_strm0 [0:4095];
  reg [31:0] pe16_lane12_strm0_tmp     ;
  reg [31:0] pe16_lane12_strm1 [0:4095];
  reg [31:0] pe16_lane12_strm1_tmp     ;
  reg [31:0] pe16_lane13_strm0 [0:4095];
  reg [31:0] pe16_lane13_strm0_tmp     ;
  reg [31:0] pe16_lane13_strm1 [0:4095];
  reg [31:0] pe16_lane13_strm1_tmp     ;
  reg [31:0] pe16_lane14_strm0 [0:4095];
  reg [31:0] pe16_lane14_strm0_tmp     ;
  reg [31:0] pe16_lane14_strm1 [0:4095];
  reg [31:0] pe16_lane14_strm1_tmp     ;
  reg [31:0] pe16_lane15_strm0 [0:4095];
  reg [31:0] pe16_lane15_strm0_tmp     ;
  reg [31:0] pe16_lane15_strm1 [0:4095];
  reg [31:0] pe16_lane15_strm1_tmp     ;
  reg [31:0] pe16_lane16_strm0 [0:4095];
  reg [31:0] pe16_lane16_strm0_tmp     ;
  reg [31:0] pe16_lane16_strm1 [0:4095];
  reg [31:0] pe16_lane16_strm1_tmp     ;
  reg [31:0] pe16_lane17_strm0 [0:4095];
  reg [31:0] pe16_lane17_strm0_tmp     ;
  reg [31:0] pe16_lane17_strm1 [0:4095];
  reg [31:0] pe16_lane17_strm1_tmp     ;
  reg [31:0] pe16_lane18_strm0 [0:4095];
  reg [31:0] pe16_lane18_strm0_tmp     ;
  reg [31:0] pe16_lane18_strm1 [0:4095];
  reg [31:0] pe16_lane18_strm1_tmp     ;
  reg [31:0] pe16_lane19_strm0 [0:4095];
  reg [31:0] pe16_lane19_strm0_tmp     ;
  reg [31:0] pe16_lane19_strm1 [0:4095];
  reg [31:0] pe16_lane19_strm1_tmp     ;
  reg [31:0] pe16_lane20_strm0 [0:4095];
  reg [31:0] pe16_lane20_strm0_tmp     ;
  reg [31:0] pe16_lane20_strm1 [0:4095];
  reg [31:0] pe16_lane20_strm1_tmp     ;
  reg [31:0] pe16_lane21_strm0 [0:4095];
  reg [31:0] pe16_lane21_strm0_tmp     ;
  reg [31:0] pe16_lane21_strm1 [0:4095];
  reg [31:0] pe16_lane21_strm1_tmp     ;
  reg [31:0] pe16_lane22_strm0 [0:4095];
  reg [31:0] pe16_lane22_strm0_tmp     ;
  reg [31:0] pe16_lane22_strm1 [0:4095];
  reg [31:0] pe16_lane22_strm1_tmp     ;
  reg [31:0] pe16_lane23_strm0 [0:4095];
  reg [31:0] pe16_lane23_strm0_tmp     ;
  reg [31:0] pe16_lane23_strm1 [0:4095];
  reg [31:0] pe16_lane23_strm1_tmp     ;
  reg [31:0] pe16_lane24_strm0 [0:4095];
  reg [31:0] pe16_lane24_strm0_tmp     ;
  reg [31:0] pe16_lane24_strm1 [0:4095];
  reg [31:0] pe16_lane24_strm1_tmp     ;
  reg [31:0] pe16_lane25_strm0 [0:4095];
  reg [31:0] pe16_lane25_strm0_tmp     ;
  reg [31:0] pe16_lane25_strm1 [0:4095];
  reg [31:0] pe16_lane25_strm1_tmp     ;
  reg [31:0] pe16_lane26_strm0 [0:4095];
  reg [31:0] pe16_lane26_strm0_tmp     ;
  reg [31:0] pe16_lane26_strm1 [0:4095];
  reg [31:0] pe16_lane26_strm1_tmp     ;
  reg [31:0] pe16_lane27_strm0 [0:4095];
  reg [31:0] pe16_lane27_strm0_tmp     ;
  reg [31:0] pe16_lane27_strm1 [0:4095];
  reg [31:0] pe16_lane27_strm1_tmp     ;
  reg [31:0] pe16_lane28_strm0 [0:4095];
  reg [31:0] pe16_lane28_strm0_tmp     ;
  reg [31:0] pe16_lane28_strm1 [0:4095];
  reg [31:0] pe16_lane28_strm1_tmp     ;
  reg [31:0] pe16_lane29_strm0 [0:4095];
  reg [31:0] pe16_lane29_strm0_tmp     ;
  reg [31:0] pe16_lane29_strm1 [0:4095];
  reg [31:0] pe16_lane29_strm1_tmp     ;
  reg [31:0] pe16_lane30_strm0 [0:4095];
  reg [31:0] pe16_lane30_strm0_tmp     ;
  reg [31:0] pe16_lane30_strm1 [0:4095];
  reg [31:0] pe16_lane30_strm1_tmp     ;
  reg [31:0] pe16_lane31_strm0 [0:4095];
  reg [31:0] pe16_lane31_strm0_tmp     ;
  reg [31:0] pe16_lane31_strm1 [0:4095];
  reg [31:0] pe16_lane31_strm1_tmp     ;
  reg [31:0] pe17_lane0_strm0 [0:4095];
  reg [31:0] pe17_lane0_strm0_tmp     ;
  reg [31:0] pe17_lane0_strm1 [0:4095];
  reg [31:0] pe17_lane0_strm1_tmp     ;
  reg [31:0] pe17_lane1_strm0 [0:4095];
  reg [31:0] pe17_lane1_strm0_tmp     ;
  reg [31:0] pe17_lane1_strm1 [0:4095];
  reg [31:0] pe17_lane1_strm1_tmp     ;
  reg [31:0] pe17_lane2_strm0 [0:4095];
  reg [31:0] pe17_lane2_strm0_tmp     ;
  reg [31:0] pe17_lane2_strm1 [0:4095];
  reg [31:0] pe17_lane2_strm1_tmp     ;
  reg [31:0] pe17_lane3_strm0 [0:4095];
  reg [31:0] pe17_lane3_strm0_tmp     ;
  reg [31:0] pe17_lane3_strm1 [0:4095];
  reg [31:0] pe17_lane3_strm1_tmp     ;
  reg [31:0] pe17_lane4_strm0 [0:4095];
  reg [31:0] pe17_lane4_strm0_tmp     ;
  reg [31:0] pe17_lane4_strm1 [0:4095];
  reg [31:0] pe17_lane4_strm1_tmp     ;
  reg [31:0] pe17_lane5_strm0 [0:4095];
  reg [31:0] pe17_lane5_strm0_tmp     ;
  reg [31:0] pe17_lane5_strm1 [0:4095];
  reg [31:0] pe17_lane5_strm1_tmp     ;
  reg [31:0] pe17_lane6_strm0 [0:4095];
  reg [31:0] pe17_lane6_strm0_tmp     ;
  reg [31:0] pe17_lane6_strm1 [0:4095];
  reg [31:0] pe17_lane6_strm1_tmp     ;
  reg [31:0] pe17_lane7_strm0 [0:4095];
  reg [31:0] pe17_lane7_strm0_tmp     ;
  reg [31:0] pe17_lane7_strm1 [0:4095];
  reg [31:0] pe17_lane7_strm1_tmp     ;
  reg [31:0] pe17_lane8_strm0 [0:4095];
  reg [31:0] pe17_lane8_strm0_tmp     ;
  reg [31:0] pe17_lane8_strm1 [0:4095];
  reg [31:0] pe17_lane8_strm1_tmp     ;
  reg [31:0] pe17_lane9_strm0 [0:4095];
  reg [31:0] pe17_lane9_strm0_tmp     ;
  reg [31:0] pe17_lane9_strm1 [0:4095];
  reg [31:0] pe17_lane9_strm1_tmp     ;
  reg [31:0] pe17_lane10_strm0 [0:4095];
  reg [31:0] pe17_lane10_strm0_tmp     ;
  reg [31:0] pe17_lane10_strm1 [0:4095];
  reg [31:0] pe17_lane10_strm1_tmp     ;
  reg [31:0] pe17_lane11_strm0 [0:4095];
  reg [31:0] pe17_lane11_strm0_tmp     ;
  reg [31:0] pe17_lane11_strm1 [0:4095];
  reg [31:0] pe17_lane11_strm1_tmp     ;
  reg [31:0] pe17_lane12_strm0 [0:4095];
  reg [31:0] pe17_lane12_strm0_tmp     ;
  reg [31:0] pe17_lane12_strm1 [0:4095];
  reg [31:0] pe17_lane12_strm1_tmp     ;
  reg [31:0] pe17_lane13_strm0 [0:4095];
  reg [31:0] pe17_lane13_strm0_tmp     ;
  reg [31:0] pe17_lane13_strm1 [0:4095];
  reg [31:0] pe17_lane13_strm1_tmp     ;
  reg [31:0] pe17_lane14_strm0 [0:4095];
  reg [31:0] pe17_lane14_strm0_tmp     ;
  reg [31:0] pe17_lane14_strm1 [0:4095];
  reg [31:0] pe17_lane14_strm1_tmp     ;
  reg [31:0] pe17_lane15_strm0 [0:4095];
  reg [31:0] pe17_lane15_strm0_tmp     ;
  reg [31:0] pe17_lane15_strm1 [0:4095];
  reg [31:0] pe17_lane15_strm1_tmp     ;
  reg [31:0] pe17_lane16_strm0 [0:4095];
  reg [31:0] pe17_lane16_strm0_tmp     ;
  reg [31:0] pe17_lane16_strm1 [0:4095];
  reg [31:0] pe17_lane16_strm1_tmp     ;
  reg [31:0] pe17_lane17_strm0 [0:4095];
  reg [31:0] pe17_lane17_strm0_tmp     ;
  reg [31:0] pe17_lane17_strm1 [0:4095];
  reg [31:0] pe17_lane17_strm1_tmp     ;
  reg [31:0] pe17_lane18_strm0 [0:4095];
  reg [31:0] pe17_lane18_strm0_tmp     ;
  reg [31:0] pe17_lane18_strm1 [0:4095];
  reg [31:0] pe17_lane18_strm1_tmp     ;
  reg [31:0] pe17_lane19_strm0 [0:4095];
  reg [31:0] pe17_lane19_strm0_tmp     ;
  reg [31:0] pe17_lane19_strm1 [0:4095];
  reg [31:0] pe17_lane19_strm1_tmp     ;
  reg [31:0] pe17_lane20_strm0 [0:4095];
  reg [31:0] pe17_lane20_strm0_tmp     ;
  reg [31:0] pe17_lane20_strm1 [0:4095];
  reg [31:0] pe17_lane20_strm1_tmp     ;
  reg [31:0] pe17_lane21_strm0 [0:4095];
  reg [31:0] pe17_lane21_strm0_tmp     ;
  reg [31:0] pe17_lane21_strm1 [0:4095];
  reg [31:0] pe17_lane21_strm1_tmp     ;
  reg [31:0] pe17_lane22_strm0 [0:4095];
  reg [31:0] pe17_lane22_strm0_tmp     ;
  reg [31:0] pe17_lane22_strm1 [0:4095];
  reg [31:0] pe17_lane22_strm1_tmp     ;
  reg [31:0] pe17_lane23_strm0 [0:4095];
  reg [31:0] pe17_lane23_strm0_tmp     ;
  reg [31:0] pe17_lane23_strm1 [0:4095];
  reg [31:0] pe17_lane23_strm1_tmp     ;
  reg [31:0] pe17_lane24_strm0 [0:4095];
  reg [31:0] pe17_lane24_strm0_tmp     ;
  reg [31:0] pe17_lane24_strm1 [0:4095];
  reg [31:0] pe17_lane24_strm1_tmp     ;
  reg [31:0] pe17_lane25_strm0 [0:4095];
  reg [31:0] pe17_lane25_strm0_tmp     ;
  reg [31:0] pe17_lane25_strm1 [0:4095];
  reg [31:0] pe17_lane25_strm1_tmp     ;
  reg [31:0] pe17_lane26_strm0 [0:4095];
  reg [31:0] pe17_lane26_strm0_tmp     ;
  reg [31:0] pe17_lane26_strm1 [0:4095];
  reg [31:0] pe17_lane26_strm1_tmp     ;
  reg [31:0] pe17_lane27_strm0 [0:4095];
  reg [31:0] pe17_lane27_strm0_tmp     ;
  reg [31:0] pe17_lane27_strm1 [0:4095];
  reg [31:0] pe17_lane27_strm1_tmp     ;
  reg [31:0] pe17_lane28_strm0 [0:4095];
  reg [31:0] pe17_lane28_strm0_tmp     ;
  reg [31:0] pe17_lane28_strm1 [0:4095];
  reg [31:0] pe17_lane28_strm1_tmp     ;
  reg [31:0] pe17_lane29_strm0 [0:4095];
  reg [31:0] pe17_lane29_strm0_tmp     ;
  reg [31:0] pe17_lane29_strm1 [0:4095];
  reg [31:0] pe17_lane29_strm1_tmp     ;
  reg [31:0] pe17_lane30_strm0 [0:4095];
  reg [31:0] pe17_lane30_strm0_tmp     ;
  reg [31:0] pe17_lane30_strm1 [0:4095];
  reg [31:0] pe17_lane30_strm1_tmp     ;
  reg [31:0] pe17_lane31_strm0 [0:4095];
  reg [31:0] pe17_lane31_strm0_tmp     ;
  reg [31:0] pe17_lane31_strm1 [0:4095];
  reg [31:0] pe17_lane31_strm1_tmp     ;
  reg [31:0] pe18_lane0_strm0 [0:4095];
  reg [31:0] pe18_lane0_strm0_tmp     ;
  reg [31:0] pe18_lane0_strm1 [0:4095];
  reg [31:0] pe18_lane0_strm1_tmp     ;
  reg [31:0] pe18_lane1_strm0 [0:4095];
  reg [31:0] pe18_lane1_strm0_tmp     ;
  reg [31:0] pe18_lane1_strm1 [0:4095];
  reg [31:0] pe18_lane1_strm1_tmp     ;
  reg [31:0] pe18_lane2_strm0 [0:4095];
  reg [31:0] pe18_lane2_strm0_tmp     ;
  reg [31:0] pe18_lane2_strm1 [0:4095];
  reg [31:0] pe18_lane2_strm1_tmp     ;
  reg [31:0] pe18_lane3_strm0 [0:4095];
  reg [31:0] pe18_lane3_strm0_tmp     ;
  reg [31:0] pe18_lane3_strm1 [0:4095];
  reg [31:0] pe18_lane3_strm1_tmp     ;
  reg [31:0] pe18_lane4_strm0 [0:4095];
  reg [31:0] pe18_lane4_strm0_tmp     ;
  reg [31:0] pe18_lane4_strm1 [0:4095];
  reg [31:0] pe18_lane4_strm1_tmp     ;
  reg [31:0] pe18_lane5_strm0 [0:4095];
  reg [31:0] pe18_lane5_strm0_tmp     ;
  reg [31:0] pe18_lane5_strm1 [0:4095];
  reg [31:0] pe18_lane5_strm1_tmp     ;
  reg [31:0] pe18_lane6_strm0 [0:4095];
  reg [31:0] pe18_lane6_strm0_tmp     ;
  reg [31:0] pe18_lane6_strm1 [0:4095];
  reg [31:0] pe18_lane6_strm1_tmp     ;
  reg [31:0] pe18_lane7_strm0 [0:4095];
  reg [31:0] pe18_lane7_strm0_tmp     ;
  reg [31:0] pe18_lane7_strm1 [0:4095];
  reg [31:0] pe18_lane7_strm1_tmp     ;
  reg [31:0] pe18_lane8_strm0 [0:4095];
  reg [31:0] pe18_lane8_strm0_tmp     ;
  reg [31:0] pe18_lane8_strm1 [0:4095];
  reg [31:0] pe18_lane8_strm1_tmp     ;
  reg [31:0] pe18_lane9_strm0 [0:4095];
  reg [31:0] pe18_lane9_strm0_tmp     ;
  reg [31:0] pe18_lane9_strm1 [0:4095];
  reg [31:0] pe18_lane9_strm1_tmp     ;
  reg [31:0] pe18_lane10_strm0 [0:4095];
  reg [31:0] pe18_lane10_strm0_tmp     ;
  reg [31:0] pe18_lane10_strm1 [0:4095];
  reg [31:0] pe18_lane10_strm1_tmp     ;
  reg [31:0] pe18_lane11_strm0 [0:4095];
  reg [31:0] pe18_lane11_strm0_tmp     ;
  reg [31:0] pe18_lane11_strm1 [0:4095];
  reg [31:0] pe18_lane11_strm1_tmp     ;
  reg [31:0] pe18_lane12_strm0 [0:4095];
  reg [31:0] pe18_lane12_strm0_tmp     ;
  reg [31:0] pe18_lane12_strm1 [0:4095];
  reg [31:0] pe18_lane12_strm1_tmp     ;
  reg [31:0] pe18_lane13_strm0 [0:4095];
  reg [31:0] pe18_lane13_strm0_tmp     ;
  reg [31:0] pe18_lane13_strm1 [0:4095];
  reg [31:0] pe18_lane13_strm1_tmp     ;
  reg [31:0] pe18_lane14_strm0 [0:4095];
  reg [31:0] pe18_lane14_strm0_tmp     ;
  reg [31:0] pe18_lane14_strm1 [0:4095];
  reg [31:0] pe18_lane14_strm1_tmp     ;
  reg [31:0] pe18_lane15_strm0 [0:4095];
  reg [31:0] pe18_lane15_strm0_tmp     ;
  reg [31:0] pe18_lane15_strm1 [0:4095];
  reg [31:0] pe18_lane15_strm1_tmp     ;
  reg [31:0] pe18_lane16_strm0 [0:4095];
  reg [31:0] pe18_lane16_strm0_tmp     ;
  reg [31:0] pe18_lane16_strm1 [0:4095];
  reg [31:0] pe18_lane16_strm1_tmp     ;
  reg [31:0] pe18_lane17_strm0 [0:4095];
  reg [31:0] pe18_lane17_strm0_tmp     ;
  reg [31:0] pe18_lane17_strm1 [0:4095];
  reg [31:0] pe18_lane17_strm1_tmp     ;
  reg [31:0] pe18_lane18_strm0 [0:4095];
  reg [31:0] pe18_lane18_strm0_tmp     ;
  reg [31:0] pe18_lane18_strm1 [0:4095];
  reg [31:0] pe18_lane18_strm1_tmp     ;
  reg [31:0] pe18_lane19_strm0 [0:4095];
  reg [31:0] pe18_lane19_strm0_tmp     ;
  reg [31:0] pe18_lane19_strm1 [0:4095];
  reg [31:0] pe18_lane19_strm1_tmp     ;
  reg [31:0] pe18_lane20_strm0 [0:4095];
  reg [31:0] pe18_lane20_strm0_tmp     ;
  reg [31:0] pe18_lane20_strm1 [0:4095];
  reg [31:0] pe18_lane20_strm1_tmp     ;
  reg [31:0] pe18_lane21_strm0 [0:4095];
  reg [31:0] pe18_lane21_strm0_tmp     ;
  reg [31:0] pe18_lane21_strm1 [0:4095];
  reg [31:0] pe18_lane21_strm1_tmp     ;
  reg [31:0] pe18_lane22_strm0 [0:4095];
  reg [31:0] pe18_lane22_strm0_tmp     ;
  reg [31:0] pe18_lane22_strm1 [0:4095];
  reg [31:0] pe18_lane22_strm1_tmp     ;
  reg [31:0] pe18_lane23_strm0 [0:4095];
  reg [31:0] pe18_lane23_strm0_tmp     ;
  reg [31:0] pe18_lane23_strm1 [0:4095];
  reg [31:0] pe18_lane23_strm1_tmp     ;
  reg [31:0] pe18_lane24_strm0 [0:4095];
  reg [31:0] pe18_lane24_strm0_tmp     ;
  reg [31:0] pe18_lane24_strm1 [0:4095];
  reg [31:0] pe18_lane24_strm1_tmp     ;
  reg [31:0] pe18_lane25_strm0 [0:4095];
  reg [31:0] pe18_lane25_strm0_tmp     ;
  reg [31:0] pe18_lane25_strm1 [0:4095];
  reg [31:0] pe18_lane25_strm1_tmp     ;
  reg [31:0] pe18_lane26_strm0 [0:4095];
  reg [31:0] pe18_lane26_strm0_tmp     ;
  reg [31:0] pe18_lane26_strm1 [0:4095];
  reg [31:0] pe18_lane26_strm1_tmp     ;
  reg [31:0] pe18_lane27_strm0 [0:4095];
  reg [31:0] pe18_lane27_strm0_tmp     ;
  reg [31:0] pe18_lane27_strm1 [0:4095];
  reg [31:0] pe18_lane27_strm1_tmp     ;
  reg [31:0] pe18_lane28_strm0 [0:4095];
  reg [31:0] pe18_lane28_strm0_tmp     ;
  reg [31:0] pe18_lane28_strm1 [0:4095];
  reg [31:0] pe18_lane28_strm1_tmp     ;
  reg [31:0] pe18_lane29_strm0 [0:4095];
  reg [31:0] pe18_lane29_strm0_tmp     ;
  reg [31:0] pe18_lane29_strm1 [0:4095];
  reg [31:0] pe18_lane29_strm1_tmp     ;
  reg [31:0] pe18_lane30_strm0 [0:4095];
  reg [31:0] pe18_lane30_strm0_tmp     ;
  reg [31:0] pe18_lane30_strm1 [0:4095];
  reg [31:0] pe18_lane30_strm1_tmp     ;
  reg [31:0] pe18_lane31_strm0 [0:4095];
  reg [31:0] pe18_lane31_strm0_tmp     ;
  reg [31:0] pe18_lane31_strm1 [0:4095];
  reg [31:0] pe18_lane31_strm1_tmp     ;
  reg [31:0] pe19_lane0_strm0 [0:4095];
  reg [31:0] pe19_lane0_strm0_tmp     ;
  reg [31:0] pe19_lane0_strm1 [0:4095];
  reg [31:0] pe19_lane0_strm1_tmp     ;
  reg [31:0] pe19_lane1_strm0 [0:4095];
  reg [31:0] pe19_lane1_strm0_tmp     ;
  reg [31:0] pe19_lane1_strm1 [0:4095];
  reg [31:0] pe19_lane1_strm1_tmp     ;
  reg [31:0] pe19_lane2_strm0 [0:4095];
  reg [31:0] pe19_lane2_strm0_tmp     ;
  reg [31:0] pe19_lane2_strm1 [0:4095];
  reg [31:0] pe19_lane2_strm1_tmp     ;
  reg [31:0] pe19_lane3_strm0 [0:4095];
  reg [31:0] pe19_lane3_strm0_tmp     ;
  reg [31:0] pe19_lane3_strm1 [0:4095];
  reg [31:0] pe19_lane3_strm1_tmp     ;
  reg [31:0] pe19_lane4_strm0 [0:4095];
  reg [31:0] pe19_lane4_strm0_tmp     ;
  reg [31:0] pe19_lane4_strm1 [0:4095];
  reg [31:0] pe19_lane4_strm1_tmp     ;
  reg [31:0] pe19_lane5_strm0 [0:4095];
  reg [31:0] pe19_lane5_strm0_tmp     ;
  reg [31:0] pe19_lane5_strm1 [0:4095];
  reg [31:0] pe19_lane5_strm1_tmp     ;
  reg [31:0] pe19_lane6_strm0 [0:4095];
  reg [31:0] pe19_lane6_strm0_tmp     ;
  reg [31:0] pe19_lane6_strm1 [0:4095];
  reg [31:0] pe19_lane6_strm1_tmp     ;
  reg [31:0] pe19_lane7_strm0 [0:4095];
  reg [31:0] pe19_lane7_strm0_tmp     ;
  reg [31:0] pe19_lane7_strm1 [0:4095];
  reg [31:0] pe19_lane7_strm1_tmp     ;
  reg [31:0] pe19_lane8_strm0 [0:4095];
  reg [31:0] pe19_lane8_strm0_tmp     ;
  reg [31:0] pe19_lane8_strm1 [0:4095];
  reg [31:0] pe19_lane8_strm1_tmp     ;
  reg [31:0] pe19_lane9_strm0 [0:4095];
  reg [31:0] pe19_lane9_strm0_tmp     ;
  reg [31:0] pe19_lane9_strm1 [0:4095];
  reg [31:0] pe19_lane9_strm1_tmp     ;
  reg [31:0] pe19_lane10_strm0 [0:4095];
  reg [31:0] pe19_lane10_strm0_tmp     ;
  reg [31:0] pe19_lane10_strm1 [0:4095];
  reg [31:0] pe19_lane10_strm1_tmp     ;
  reg [31:0] pe19_lane11_strm0 [0:4095];
  reg [31:0] pe19_lane11_strm0_tmp     ;
  reg [31:0] pe19_lane11_strm1 [0:4095];
  reg [31:0] pe19_lane11_strm1_tmp     ;
  reg [31:0] pe19_lane12_strm0 [0:4095];
  reg [31:0] pe19_lane12_strm0_tmp     ;
  reg [31:0] pe19_lane12_strm1 [0:4095];
  reg [31:0] pe19_lane12_strm1_tmp     ;
  reg [31:0] pe19_lane13_strm0 [0:4095];
  reg [31:0] pe19_lane13_strm0_tmp     ;
  reg [31:0] pe19_lane13_strm1 [0:4095];
  reg [31:0] pe19_lane13_strm1_tmp     ;
  reg [31:0] pe19_lane14_strm0 [0:4095];
  reg [31:0] pe19_lane14_strm0_tmp     ;
  reg [31:0] pe19_lane14_strm1 [0:4095];
  reg [31:0] pe19_lane14_strm1_tmp     ;
  reg [31:0] pe19_lane15_strm0 [0:4095];
  reg [31:0] pe19_lane15_strm0_tmp     ;
  reg [31:0] pe19_lane15_strm1 [0:4095];
  reg [31:0] pe19_lane15_strm1_tmp     ;
  reg [31:0] pe19_lane16_strm0 [0:4095];
  reg [31:0] pe19_lane16_strm0_tmp     ;
  reg [31:0] pe19_lane16_strm1 [0:4095];
  reg [31:0] pe19_lane16_strm1_tmp     ;
  reg [31:0] pe19_lane17_strm0 [0:4095];
  reg [31:0] pe19_lane17_strm0_tmp     ;
  reg [31:0] pe19_lane17_strm1 [0:4095];
  reg [31:0] pe19_lane17_strm1_tmp     ;
  reg [31:0] pe19_lane18_strm0 [0:4095];
  reg [31:0] pe19_lane18_strm0_tmp     ;
  reg [31:0] pe19_lane18_strm1 [0:4095];
  reg [31:0] pe19_lane18_strm1_tmp     ;
  reg [31:0] pe19_lane19_strm0 [0:4095];
  reg [31:0] pe19_lane19_strm0_tmp     ;
  reg [31:0] pe19_lane19_strm1 [0:4095];
  reg [31:0] pe19_lane19_strm1_tmp     ;
  reg [31:0] pe19_lane20_strm0 [0:4095];
  reg [31:0] pe19_lane20_strm0_tmp     ;
  reg [31:0] pe19_lane20_strm1 [0:4095];
  reg [31:0] pe19_lane20_strm1_tmp     ;
  reg [31:0] pe19_lane21_strm0 [0:4095];
  reg [31:0] pe19_lane21_strm0_tmp     ;
  reg [31:0] pe19_lane21_strm1 [0:4095];
  reg [31:0] pe19_lane21_strm1_tmp     ;
  reg [31:0] pe19_lane22_strm0 [0:4095];
  reg [31:0] pe19_lane22_strm0_tmp     ;
  reg [31:0] pe19_lane22_strm1 [0:4095];
  reg [31:0] pe19_lane22_strm1_tmp     ;
  reg [31:0] pe19_lane23_strm0 [0:4095];
  reg [31:0] pe19_lane23_strm0_tmp     ;
  reg [31:0] pe19_lane23_strm1 [0:4095];
  reg [31:0] pe19_lane23_strm1_tmp     ;
  reg [31:0] pe19_lane24_strm0 [0:4095];
  reg [31:0] pe19_lane24_strm0_tmp     ;
  reg [31:0] pe19_lane24_strm1 [0:4095];
  reg [31:0] pe19_lane24_strm1_tmp     ;
  reg [31:0] pe19_lane25_strm0 [0:4095];
  reg [31:0] pe19_lane25_strm0_tmp     ;
  reg [31:0] pe19_lane25_strm1 [0:4095];
  reg [31:0] pe19_lane25_strm1_tmp     ;
  reg [31:0] pe19_lane26_strm0 [0:4095];
  reg [31:0] pe19_lane26_strm0_tmp     ;
  reg [31:0] pe19_lane26_strm1 [0:4095];
  reg [31:0] pe19_lane26_strm1_tmp     ;
  reg [31:0] pe19_lane27_strm0 [0:4095];
  reg [31:0] pe19_lane27_strm0_tmp     ;
  reg [31:0] pe19_lane27_strm1 [0:4095];
  reg [31:0] pe19_lane27_strm1_tmp     ;
  reg [31:0] pe19_lane28_strm0 [0:4095];
  reg [31:0] pe19_lane28_strm0_tmp     ;
  reg [31:0] pe19_lane28_strm1 [0:4095];
  reg [31:0] pe19_lane28_strm1_tmp     ;
  reg [31:0] pe19_lane29_strm0 [0:4095];
  reg [31:0] pe19_lane29_strm0_tmp     ;
  reg [31:0] pe19_lane29_strm1 [0:4095];
  reg [31:0] pe19_lane29_strm1_tmp     ;
  reg [31:0] pe19_lane30_strm0 [0:4095];
  reg [31:0] pe19_lane30_strm0_tmp     ;
  reg [31:0] pe19_lane30_strm1 [0:4095];
  reg [31:0] pe19_lane30_strm1_tmp     ;
  reg [31:0] pe19_lane31_strm0 [0:4095];
  reg [31:0] pe19_lane31_strm0_tmp     ;
  reg [31:0] pe19_lane31_strm1 [0:4095];
  reg [31:0] pe19_lane31_strm1_tmp     ;
  reg [31:0] pe20_lane0_strm0 [0:4095];
  reg [31:0] pe20_lane0_strm0_tmp     ;
  reg [31:0] pe20_lane0_strm1 [0:4095];
  reg [31:0] pe20_lane0_strm1_tmp     ;
  reg [31:0] pe20_lane1_strm0 [0:4095];
  reg [31:0] pe20_lane1_strm0_tmp     ;
  reg [31:0] pe20_lane1_strm1 [0:4095];
  reg [31:0] pe20_lane1_strm1_tmp     ;
  reg [31:0] pe20_lane2_strm0 [0:4095];
  reg [31:0] pe20_lane2_strm0_tmp     ;
  reg [31:0] pe20_lane2_strm1 [0:4095];
  reg [31:0] pe20_lane2_strm1_tmp     ;
  reg [31:0] pe20_lane3_strm0 [0:4095];
  reg [31:0] pe20_lane3_strm0_tmp     ;
  reg [31:0] pe20_lane3_strm1 [0:4095];
  reg [31:0] pe20_lane3_strm1_tmp     ;
  reg [31:0] pe20_lane4_strm0 [0:4095];
  reg [31:0] pe20_lane4_strm0_tmp     ;
  reg [31:0] pe20_lane4_strm1 [0:4095];
  reg [31:0] pe20_lane4_strm1_tmp     ;
  reg [31:0] pe20_lane5_strm0 [0:4095];
  reg [31:0] pe20_lane5_strm0_tmp     ;
  reg [31:0] pe20_lane5_strm1 [0:4095];
  reg [31:0] pe20_lane5_strm1_tmp     ;
  reg [31:0] pe20_lane6_strm0 [0:4095];
  reg [31:0] pe20_lane6_strm0_tmp     ;
  reg [31:0] pe20_lane6_strm1 [0:4095];
  reg [31:0] pe20_lane6_strm1_tmp     ;
  reg [31:0] pe20_lane7_strm0 [0:4095];
  reg [31:0] pe20_lane7_strm0_tmp     ;
  reg [31:0] pe20_lane7_strm1 [0:4095];
  reg [31:0] pe20_lane7_strm1_tmp     ;
  reg [31:0] pe20_lane8_strm0 [0:4095];
  reg [31:0] pe20_lane8_strm0_tmp     ;
  reg [31:0] pe20_lane8_strm1 [0:4095];
  reg [31:0] pe20_lane8_strm1_tmp     ;
  reg [31:0] pe20_lane9_strm0 [0:4095];
  reg [31:0] pe20_lane9_strm0_tmp     ;
  reg [31:0] pe20_lane9_strm1 [0:4095];
  reg [31:0] pe20_lane9_strm1_tmp     ;
  reg [31:0] pe20_lane10_strm0 [0:4095];
  reg [31:0] pe20_lane10_strm0_tmp     ;
  reg [31:0] pe20_lane10_strm1 [0:4095];
  reg [31:0] pe20_lane10_strm1_tmp     ;
  reg [31:0] pe20_lane11_strm0 [0:4095];
  reg [31:0] pe20_lane11_strm0_tmp     ;
  reg [31:0] pe20_lane11_strm1 [0:4095];
  reg [31:0] pe20_lane11_strm1_tmp     ;
  reg [31:0] pe20_lane12_strm0 [0:4095];
  reg [31:0] pe20_lane12_strm0_tmp     ;
  reg [31:0] pe20_lane12_strm1 [0:4095];
  reg [31:0] pe20_lane12_strm1_tmp     ;
  reg [31:0] pe20_lane13_strm0 [0:4095];
  reg [31:0] pe20_lane13_strm0_tmp     ;
  reg [31:0] pe20_lane13_strm1 [0:4095];
  reg [31:0] pe20_lane13_strm1_tmp     ;
  reg [31:0] pe20_lane14_strm0 [0:4095];
  reg [31:0] pe20_lane14_strm0_tmp     ;
  reg [31:0] pe20_lane14_strm1 [0:4095];
  reg [31:0] pe20_lane14_strm1_tmp     ;
  reg [31:0] pe20_lane15_strm0 [0:4095];
  reg [31:0] pe20_lane15_strm0_tmp     ;
  reg [31:0] pe20_lane15_strm1 [0:4095];
  reg [31:0] pe20_lane15_strm1_tmp     ;
  reg [31:0] pe20_lane16_strm0 [0:4095];
  reg [31:0] pe20_lane16_strm0_tmp     ;
  reg [31:0] pe20_lane16_strm1 [0:4095];
  reg [31:0] pe20_lane16_strm1_tmp     ;
  reg [31:0] pe20_lane17_strm0 [0:4095];
  reg [31:0] pe20_lane17_strm0_tmp     ;
  reg [31:0] pe20_lane17_strm1 [0:4095];
  reg [31:0] pe20_lane17_strm1_tmp     ;
  reg [31:0] pe20_lane18_strm0 [0:4095];
  reg [31:0] pe20_lane18_strm0_tmp     ;
  reg [31:0] pe20_lane18_strm1 [0:4095];
  reg [31:0] pe20_lane18_strm1_tmp     ;
  reg [31:0] pe20_lane19_strm0 [0:4095];
  reg [31:0] pe20_lane19_strm0_tmp     ;
  reg [31:0] pe20_lane19_strm1 [0:4095];
  reg [31:0] pe20_lane19_strm1_tmp     ;
  reg [31:0] pe20_lane20_strm0 [0:4095];
  reg [31:0] pe20_lane20_strm0_tmp     ;
  reg [31:0] pe20_lane20_strm1 [0:4095];
  reg [31:0] pe20_lane20_strm1_tmp     ;
  reg [31:0] pe20_lane21_strm0 [0:4095];
  reg [31:0] pe20_lane21_strm0_tmp     ;
  reg [31:0] pe20_lane21_strm1 [0:4095];
  reg [31:0] pe20_lane21_strm1_tmp     ;
  reg [31:0] pe20_lane22_strm0 [0:4095];
  reg [31:0] pe20_lane22_strm0_tmp     ;
  reg [31:0] pe20_lane22_strm1 [0:4095];
  reg [31:0] pe20_lane22_strm1_tmp     ;
  reg [31:0] pe20_lane23_strm0 [0:4095];
  reg [31:0] pe20_lane23_strm0_tmp     ;
  reg [31:0] pe20_lane23_strm1 [0:4095];
  reg [31:0] pe20_lane23_strm1_tmp     ;
  reg [31:0] pe20_lane24_strm0 [0:4095];
  reg [31:0] pe20_lane24_strm0_tmp     ;
  reg [31:0] pe20_lane24_strm1 [0:4095];
  reg [31:0] pe20_lane24_strm1_tmp     ;
  reg [31:0] pe20_lane25_strm0 [0:4095];
  reg [31:0] pe20_lane25_strm0_tmp     ;
  reg [31:0] pe20_lane25_strm1 [0:4095];
  reg [31:0] pe20_lane25_strm1_tmp     ;
  reg [31:0] pe20_lane26_strm0 [0:4095];
  reg [31:0] pe20_lane26_strm0_tmp     ;
  reg [31:0] pe20_lane26_strm1 [0:4095];
  reg [31:0] pe20_lane26_strm1_tmp     ;
  reg [31:0] pe20_lane27_strm0 [0:4095];
  reg [31:0] pe20_lane27_strm0_tmp     ;
  reg [31:0] pe20_lane27_strm1 [0:4095];
  reg [31:0] pe20_lane27_strm1_tmp     ;
  reg [31:0] pe20_lane28_strm0 [0:4095];
  reg [31:0] pe20_lane28_strm0_tmp     ;
  reg [31:0] pe20_lane28_strm1 [0:4095];
  reg [31:0] pe20_lane28_strm1_tmp     ;
  reg [31:0] pe20_lane29_strm0 [0:4095];
  reg [31:0] pe20_lane29_strm0_tmp     ;
  reg [31:0] pe20_lane29_strm1 [0:4095];
  reg [31:0] pe20_lane29_strm1_tmp     ;
  reg [31:0] pe20_lane30_strm0 [0:4095];
  reg [31:0] pe20_lane30_strm0_tmp     ;
  reg [31:0] pe20_lane30_strm1 [0:4095];
  reg [31:0] pe20_lane30_strm1_tmp     ;
  reg [31:0] pe20_lane31_strm0 [0:4095];
  reg [31:0] pe20_lane31_strm0_tmp     ;
  reg [31:0] pe20_lane31_strm1 [0:4095];
  reg [31:0] pe20_lane31_strm1_tmp     ;
  reg [31:0] pe21_lane0_strm0 [0:4095];
  reg [31:0] pe21_lane0_strm0_tmp     ;
  reg [31:0] pe21_lane0_strm1 [0:4095];
  reg [31:0] pe21_lane0_strm1_tmp     ;
  reg [31:0] pe21_lane1_strm0 [0:4095];
  reg [31:0] pe21_lane1_strm0_tmp     ;
  reg [31:0] pe21_lane1_strm1 [0:4095];
  reg [31:0] pe21_lane1_strm1_tmp     ;
  reg [31:0] pe21_lane2_strm0 [0:4095];
  reg [31:0] pe21_lane2_strm0_tmp     ;
  reg [31:0] pe21_lane2_strm1 [0:4095];
  reg [31:0] pe21_lane2_strm1_tmp     ;
  reg [31:0] pe21_lane3_strm0 [0:4095];
  reg [31:0] pe21_lane3_strm0_tmp     ;
  reg [31:0] pe21_lane3_strm1 [0:4095];
  reg [31:0] pe21_lane3_strm1_tmp     ;
  reg [31:0] pe21_lane4_strm0 [0:4095];
  reg [31:0] pe21_lane4_strm0_tmp     ;
  reg [31:0] pe21_lane4_strm1 [0:4095];
  reg [31:0] pe21_lane4_strm1_tmp     ;
  reg [31:0] pe21_lane5_strm0 [0:4095];
  reg [31:0] pe21_lane5_strm0_tmp     ;
  reg [31:0] pe21_lane5_strm1 [0:4095];
  reg [31:0] pe21_lane5_strm1_tmp     ;
  reg [31:0] pe21_lane6_strm0 [0:4095];
  reg [31:0] pe21_lane6_strm0_tmp     ;
  reg [31:0] pe21_lane6_strm1 [0:4095];
  reg [31:0] pe21_lane6_strm1_tmp     ;
  reg [31:0] pe21_lane7_strm0 [0:4095];
  reg [31:0] pe21_lane7_strm0_tmp     ;
  reg [31:0] pe21_lane7_strm1 [0:4095];
  reg [31:0] pe21_lane7_strm1_tmp     ;
  reg [31:0] pe21_lane8_strm0 [0:4095];
  reg [31:0] pe21_lane8_strm0_tmp     ;
  reg [31:0] pe21_lane8_strm1 [0:4095];
  reg [31:0] pe21_lane8_strm1_tmp     ;
  reg [31:0] pe21_lane9_strm0 [0:4095];
  reg [31:0] pe21_lane9_strm0_tmp     ;
  reg [31:0] pe21_lane9_strm1 [0:4095];
  reg [31:0] pe21_lane9_strm1_tmp     ;
  reg [31:0] pe21_lane10_strm0 [0:4095];
  reg [31:0] pe21_lane10_strm0_tmp     ;
  reg [31:0] pe21_lane10_strm1 [0:4095];
  reg [31:0] pe21_lane10_strm1_tmp     ;
  reg [31:0] pe21_lane11_strm0 [0:4095];
  reg [31:0] pe21_lane11_strm0_tmp     ;
  reg [31:0] pe21_lane11_strm1 [0:4095];
  reg [31:0] pe21_lane11_strm1_tmp     ;
  reg [31:0] pe21_lane12_strm0 [0:4095];
  reg [31:0] pe21_lane12_strm0_tmp     ;
  reg [31:0] pe21_lane12_strm1 [0:4095];
  reg [31:0] pe21_lane12_strm1_tmp     ;
  reg [31:0] pe21_lane13_strm0 [0:4095];
  reg [31:0] pe21_lane13_strm0_tmp     ;
  reg [31:0] pe21_lane13_strm1 [0:4095];
  reg [31:0] pe21_lane13_strm1_tmp     ;
  reg [31:0] pe21_lane14_strm0 [0:4095];
  reg [31:0] pe21_lane14_strm0_tmp     ;
  reg [31:0] pe21_lane14_strm1 [0:4095];
  reg [31:0] pe21_lane14_strm1_tmp     ;
  reg [31:0] pe21_lane15_strm0 [0:4095];
  reg [31:0] pe21_lane15_strm0_tmp     ;
  reg [31:0] pe21_lane15_strm1 [0:4095];
  reg [31:0] pe21_lane15_strm1_tmp     ;
  reg [31:0] pe21_lane16_strm0 [0:4095];
  reg [31:0] pe21_lane16_strm0_tmp     ;
  reg [31:0] pe21_lane16_strm1 [0:4095];
  reg [31:0] pe21_lane16_strm1_tmp     ;
  reg [31:0] pe21_lane17_strm0 [0:4095];
  reg [31:0] pe21_lane17_strm0_tmp     ;
  reg [31:0] pe21_lane17_strm1 [0:4095];
  reg [31:0] pe21_lane17_strm1_tmp     ;
  reg [31:0] pe21_lane18_strm0 [0:4095];
  reg [31:0] pe21_lane18_strm0_tmp     ;
  reg [31:0] pe21_lane18_strm1 [0:4095];
  reg [31:0] pe21_lane18_strm1_tmp     ;
  reg [31:0] pe21_lane19_strm0 [0:4095];
  reg [31:0] pe21_lane19_strm0_tmp     ;
  reg [31:0] pe21_lane19_strm1 [0:4095];
  reg [31:0] pe21_lane19_strm1_tmp     ;
  reg [31:0] pe21_lane20_strm0 [0:4095];
  reg [31:0] pe21_lane20_strm0_tmp     ;
  reg [31:0] pe21_lane20_strm1 [0:4095];
  reg [31:0] pe21_lane20_strm1_tmp     ;
  reg [31:0] pe21_lane21_strm0 [0:4095];
  reg [31:0] pe21_lane21_strm0_tmp     ;
  reg [31:0] pe21_lane21_strm1 [0:4095];
  reg [31:0] pe21_lane21_strm1_tmp     ;
  reg [31:0] pe21_lane22_strm0 [0:4095];
  reg [31:0] pe21_lane22_strm0_tmp     ;
  reg [31:0] pe21_lane22_strm1 [0:4095];
  reg [31:0] pe21_lane22_strm1_tmp     ;
  reg [31:0] pe21_lane23_strm0 [0:4095];
  reg [31:0] pe21_lane23_strm0_tmp     ;
  reg [31:0] pe21_lane23_strm1 [0:4095];
  reg [31:0] pe21_lane23_strm1_tmp     ;
  reg [31:0] pe21_lane24_strm0 [0:4095];
  reg [31:0] pe21_lane24_strm0_tmp     ;
  reg [31:0] pe21_lane24_strm1 [0:4095];
  reg [31:0] pe21_lane24_strm1_tmp     ;
  reg [31:0] pe21_lane25_strm0 [0:4095];
  reg [31:0] pe21_lane25_strm0_tmp     ;
  reg [31:0] pe21_lane25_strm1 [0:4095];
  reg [31:0] pe21_lane25_strm1_tmp     ;
  reg [31:0] pe21_lane26_strm0 [0:4095];
  reg [31:0] pe21_lane26_strm0_tmp     ;
  reg [31:0] pe21_lane26_strm1 [0:4095];
  reg [31:0] pe21_lane26_strm1_tmp     ;
  reg [31:0] pe21_lane27_strm0 [0:4095];
  reg [31:0] pe21_lane27_strm0_tmp     ;
  reg [31:0] pe21_lane27_strm1 [0:4095];
  reg [31:0] pe21_lane27_strm1_tmp     ;
  reg [31:0] pe21_lane28_strm0 [0:4095];
  reg [31:0] pe21_lane28_strm0_tmp     ;
  reg [31:0] pe21_lane28_strm1 [0:4095];
  reg [31:0] pe21_lane28_strm1_tmp     ;
  reg [31:0] pe21_lane29_strm0 [0:4095];
  reg [31:0] pe21_lane29_strm0_tmp     ;
  reg [31:0] pe21_lane29_strm1 [0:4095];
  reg [31:0] pe21_lane29_strm1_tmp     ;
  reg [31:0] pe21_lane30_strm0 [0:4095];
  reg [31:0] pe21_lane30_strm0_tmp     ;
  reg [31:0] pe21_lane30_strm1 [0:4095];
  reg [31:0] pe21_lane30_strm1_tmp     ;
  reg [31:0] pe21_lane31_strm0 [0:4095];
  reg [31:0] pe21_lane31_strm0_tmp     ;
  reg [31:0] pe21_lane31_strm1 [0:4095];
  reg [31:0] pe21_lane31_strm1_tmp     ;
  reg [31:0] pe22_lane0_strm0 [0:4095];
  reg [31:0] pe22_lane0_strm0_tmp     ;
  reg [31:0] pe22_lane0_strm1 [0:4095];
  reg [31:0] pe22_lane0_strm1_tmp     ;
  reg [31:0] pe22_lane1_strm0 [0:4095];
  reg [31:0] pe22_lane1_strm0_tmp     ;
  reg [31:0] pe22_lane1_strm1 [0:4095];
  reg [31:0] pe22_lane1_strm1_tmp     ;
  reg [31:0] pe22_lane2_strm0 [0:4095];
  reg [31:0] pe22_lane2_strm0_tmp     ;
  reg [31:0] pe22_lane2_strm1 [0:4095];
  reg [31:0] pe22_lane2_strm1_tmp     ;
  reg [31:0] pe22_lane3_strm0 [0:4095];
  reg [31:0] pe22_lane3_strm0_tmp     ;
  reg [31:0] pe22_lane3_strm1 [0:4095];
  reg [31:0] pe22_lane3_strm1_tmp     ;
  reg [31:0] pe22_lane4_strm0 [0:4095];
  reg [31:0] pe22_lane4_strm0_tmp     ;
  reg [31:0] pe22_lane4_strm1 [0:4095];
  reg [31:0] pe22_lane4_strm1_tmp     ;
  reg [31:0] pe22_lane5_strm0 [0:4095];
  reg [31:0] pe22_lane5_strm0_tmp     ;
  reg [31:0] pe22_lane5_strm1 [0:4095];
  reg [31:0] pe22_lane5_strm1_tmp     ;
  reg [31:0] pe22_lane6_strm0 [0:4095];
  reg [31:0] pe22_lane6_strm0_tmp     ;
  reg [31:0] pe22_lane6_strm1 [0:4095];
  reg [31:0] pe22_lane6_strm1_tmp     ;
  reg [31:0] pe22_lane7_strm0 [0:4095];
  reg [31:0] pe22_lane7_strm0_tmp     ;
  reg [31:0] pe22_lane7_strm1 [0:4095];
  reg [31:0] pe22_lane7_strm1_tmp     ;
  reg [31:0] pe22_lane8_strm0 [0:4095];
  reg [31:0] pe22_lane8_strm0_tmp     ;
  reg [31:0] pe22_lane8_strm1 [0:4095];
  reg [31:0] pe22_lane8_strm1_tmp     ;
  reg [31:0] pe22_lane9_strm0 [0:4095];
  reg [31:0] pe22_lane9_strm0_tmp     ;
  reg [31:0] pe22_lane9_strm1 [0:4095];
  reg [31:0] pe22_lane9_strm1_tmp     ;
  reg [31:0] pe22_lane10_strm0 [0:4095];
  reg [31:0] pe22_lane10_strm0_tmp     ;
  reg [31:0] pe22_lane10_strm1 [0:4095];
  reg [31:0] pe22_lane10_strm1_tmp     ;
  reg [31:0] pe22_lane11_strm0 [0:4095];
  reg [31:0] pe22_lane11_strm0_tmp     ;
  reg [31:0] pe22_lane11_strm1 [0:4095];
  reg [31:0] pe22_lane11_strm1_tmp     ;
  reg [31:0] pe22_lane12_strm0 [0:4095];
  reg [31:0] pe22_lane12_strm0_tmp     ;
  reg [31:0] pe22_lane12_strm1 [0:4095];
  reg [31:0] pe22_lane12_strm1_tmp     ;
  reg [31:0] pe22_lane13_strm0 [0:4095];
  reg [31:0] pe22_lane13_strm0_tmp     ;
  reg [31:0] pe22_lane13_strm1 [0:4095];
  reg [31:0] pe22_lane13_strm1_tmp     ;
  reg [31:0] pe22_lane14_strm0 [0:4095];
  reg [31:0] pe22_lane14_strm0_tmp     ;
  reg [31:0] pe22_lane14_strm1 [0:4095];
  reg [31:0] pe22_lane14_strm1_tmp     ;
  reg [31:0] pe22_lane15_strm0 [0:4095];
  reg [31:0] pe22_lane15_strm0_tmp     ;
  reg [31:0] pe22_lane15_strm1 [0:4095];
  reg [31:0] pe22_lane15_strm1_tmp     ;
  reg [31:0] pe22_lane16_strm0 [0:4095];
  reg [31:0] pe22_lane16_strm0_tmp     ;
  reg [31:0] pe22_lane16_strm1 [0:4095];
  reg [31:0] pe22_lane16_strm1_tmp     ;
  reg [31:0] pe22_lane17_strm0 [0:4095];
  reg [31:0] pe22_lane17_strm0_tmp     ;
  reg [31:0] pe22_lane17_strm1 [0:4095];
  reg [31:0] pe22_lane17_strm1_tmp     ;
  reg [31:0] pe22_lane18_strm0 [0:4095];
  reg [31:0] pe22_lane18_strm0_tmp     ;
  reg [31:0] pe22_lane18_strm1 [0:4095];
  reg [31:0] pe22_lane18_strm1_tmp     ;
  reg [31:0] pe22_lane19_strm0 [0:4095];
  reg [31:0] pe22_lane19_strm0_tmp     ;
  reg [31:0] pe22_lane19_strm1 [0:4095];
  reg [31:0] pe22_lane19_strm1_tmp     ;
  reg [31:0] pe22_lane20_strm0 [0:4095];
  reg [31:0] pe22_lane20_strm0_tmp     ;
  reg [31:0] pe22_lane20_strm1 [0:4095];
  reg [31:0] pe22_lane20_strm1_tmp     ;
  reg [31:0] pe22_lane21_strm0 [0:4095];
  reg [31:0] pe22_lane21_strm0_tmp     ;
  reg [31:0] pe22_lane21_strm1 [0:4095];
  reg [31:0] pe22_lane21_strm1_tmp     ;
  reg [31:0] pe22_lane22_strm0 [0:4095];
  reg [31:0] pe22_lane22_strm0_tmp     ;
  reg [31:0] pe22_lane22_strm1 [0:4095];
  reg [31:0] pe22_lane22_strm1_tmp     ;
  reg [31:0] pe22_lane23_strm0 [0:4095];
  reg [31:0] pe22_lane23_strm0_tmp     ;
  reg [31:0] pe22_lane23_strm1 [0:4095];
  reg [31:0] pe22_lane23_strm1_tmp     ;
  reg [31:0] pe22_lane24_strm0 [0:4095];
  reg [31:0] pe22_lane24_strm0_tmp     ;
  reg [31:0] pe22_lane24_strm1 [0:4095];
  reg [31:0] pe22_lane24_strm1_tmp     ;
  reg [31:0] pe22_lane25_strm0 [0:4095];
  reg [31:0] pe22_lane25_strm0_tmp     ;
  reg [31:0] pe22_lane25_strm1 [0:4095];
  reg [31:0] pe22_lane25_strm1_tmp     ;
  reg [31:0] pe22_lane26_strm0 [0:4095];
  reg [31:0] pe22_lane26_strm0_tmp     ;
  reg [31:0] pe22_lane26_strm1 [0:4095];
  reg [31:0] pe22_lane26_strm1_tmp     ;
  reg [31:0] pe22_lane27_strm0 [0:4095];
  reg [31:0] pe22_lane27_strm0_tmp     ;
  reg [31:0] pe22_lane27_strm1 [0:4095];
  reg [31:0] pe22_lane27_strm1_tmp     ;
  reg [31:0] pe22_lane28_strm0 [0:4095];
  reg [31:0] pe22_lane28_strm0_tmp     ;
  reg [31:0] pe22_lane28_strm1 [0:4095];
  reg [31:0] pe22_lane28_strm1_tmp     ;
  reg [31:0] pe22_lane29_strm0 [0:4095];
  reg [31:0] pe22_lane29_strm0_tmp     ;
  reg [31:0] pe22_lane29_strm1 [0:4095];
  reg [31:0] pe22_lane29_strm1_tmp     ;
  reg [31:0] pe22_lane30_strm0 [0:4095];
  reg [31:0] pe22_lane30_strm0_tmp     ;
  reg [31:0] pe22_lane30_strm1 [0:4095];
  reg [31:0] pe22_lane30_strm1_tmp     ;
  reg [31:0] pe22_lane31_strm0 [0:4095];
  reg [31:0] pe22_lane31_strm0_tmp     ;
  reg [31:0] pe22_lane31_strm1 [0:4095];
  reg [31:0] pe22_lane31_strm1_tmp     ;
  reg [31:0] pe23_lane0_strm0 [0:4095];
  reg [31:0] pe23_lane0_strm0_tmp     ;
  reg [31:0] pe23_lane0_strm1 [0:4095];
  reg [31:0] pe23_lane0_strm1_tmp     ;
  reg [31:0] pe23_lane1_strm0 [0:4095];
  reg [31:0] pe23_lane1_strm0_tmp     ;
  reg [31:0] pe23_lane1_strm1 [0:4095];
  reg [31:0] pe23_lane1_strm1_tmp     ;
  reg [31:0] pe23_lane2_strm0 [0:4095];
  reg [31:0] pe23_lane2_strm0_tmp     ;
  reg [31:0] pe23_lane2_strm1 [0:4095];
  reg [31:0] pe23_lane2_strm1_tmp     ;
  reg [31:0] pe23_lane3_strm0 [0:4095];
  reg [31:0] pe23_lane3_strm0_tmp     ;
  reg [31:0] pe23_lane3_strm1 [0:4095];
  reg [31:0] pe23_lane3_strm1_tmp     ;
  reg [31:0] pe23_lane4_strm0 [0:4095];
  reg [31:0] pe23_lane4_strm0_tmp     ;
  reg [31:0] pe23_lane4_strm1 [0:4095];
  reg [31:0] pe23_lane4_strm1_tmp     ;
  reg [31:0] pe23_lane5_strm0 [0:4095];
  reg [31:0] pe23_lane5_strm0_tmp     ;
  reg [31:0] pe23_lane5_strm1 [0:4095];
  reg [31:0] pe23_lane5_strm1_tmp     ;
  reg [31:0] pe23_lane6_strm0 [0:4095];
  reg [31:0] pe23_lane6_strm0_tmp     ;
  reg [31:0] pe23_lane6_strm1 [0:4095];
  reg [31:0] pe23_lane6_strm1_tmp     ;
  reg [31:0] pe23_lane7_strm0 [0:4095];
  reg [31:0] pe23_lane7_strm0_tmp     ;
  reg [31:0] pe23_lane7_strm1 [0:4095];
  reg [31:0] pe23_lane7_strm1_tmp     ;
  reg [31:0] pe23_lane8_strm0 [0:4095];
  reg [31:0] pe23_lane8_strm0_tmp     ;
  reg [31:0] pe23_lane8_strm1 [0:4095];
  reg [31:0] pe23_lane8_strm1_tmp     ;
  reg [31:0] pe23_lane9_strm0 [0:4095];
  reg [31:0] pe23_lane9_strm0_tmp     ;
  reg [31:0] pe23_lane9_strm1 [0:4095];
  reg [31:0] pe23_lane9_strm1_tmp     ;
  reg [31:0] pe23_lane10_strm0 [0:4095];
  reg [31:0] pe23_lane10_strm0_tmp     ;
  reg [31:0] pe23_lane10_strm1 [0:4095];
  reg [31:0] pe23_lane10_strm1_tmp     ;
  reg [31:0] pe23_lane11_strm0 [0:4095];
  reg [31:0] pe23_lane11_strm0_tmp     ;
  reg [31:0] pe23_lane11_strm1 [0:4095];
  reg [31:0] pe23_lane11_strm1_tmp     ;
  reg [31:0] pe23_lane12_strm0 [0:4095];
  reg [31:0] pe23_lane12_strm0_tmp     ;
  reg [31:0] pe23_lane12_strm1 [0:4095];
  reg [31:0] pe23_lane12_strm1_tmp     ;
  reg [31:0] pe23_lane13_strm0 [0:4095];
  reg [31:0] pe23_lane13_strm0_tmp     ;
  reg [31:0] pe23_lane13_strm1 [0:4095];
  reg [31:0] pe23_lane13_strm1_tmp     ;
  reg [31:0] pe23_lane14_strm0 [0:4095];
  reg [31:0] pe23_lane14_strm0_tmp     ;
  reg [31:0] pe23_lane14_strm1 [0:4095];
  reg [31:0] pe23_lane14_strm1_tmp     ;
  reg [31:0] pe23_lane15_strm0 [0:4095];
  reg [31:0] pe23_lane15_strm0_tmp     ;
  reg [31:0] pe23_lane15_strm1 [0:4095];
  reg [31:0] pe23_lane15_strm1_tmp     ;
  reg [31:0] pe23_lane16_strm0 [0:4095];
  reg [31:0] pe23_lane16_strm0_tmp     ;
  reg [31:0] pe23_lane16_strm1 [0:4095];
  reg [31:0] pe23_lane16_strm1_tmp     ;
  reg [31:0] pe23_lane17_strm0 [0:4095];
  reg [31:0] pe23_lane17_strm0_tmp     ;
  reg [31:0] pe23_lane17_strm1 [0:4095];
  reg [31:0] pe23_lane17_strm1_tmp     ;
  reg [31:0] pe23_lane18_strm0 [0:4095];
  reg [31:0] pe23_lane18_strm0_tmp     ;
  reg [31:0] pe23_lane18_strm1 [0:4095];
  reg [31:0] pe23_lane18_strm1_tmp     ;
  reg [31:0] pe23_lane19_strm0 [0:4095];
  reg [31:0] pe23_lane19_strm0_tmp     ;
  reg [31:0] pe23_lane19_strm1 [0:4095];
  reg [31:0] pe23_lane19_strm1_tmp     ;
  reg [31:0] pe23_lane20_strm0 [0:4095];
  reg [31:0] pe23_lane20_strm0_tmp     ;
  reg [31:0] pe23_lane20_strm1 [0:4095];
  reg [31:0] pe23_lane20_strm1_tmp     ;
  reg [31:0] pe23_lane21_strm0 [0:4095];
  reg [31:0] pe23_lane21_strm0_tmp     ;
  reg [31:0] pe23_lane21_strm1 [0:4095];
  reg [31:0] pe23_lane21_strm1_tmp     ;
  reg [31:0] pe23_lane22_strm0 [0:4095];
  reg [31:0] pe23_lane22_strm0_tmp     ;
  reg [31:0] pe23_lane22_strm1 [0:4095];
  reg [31:0] pe23_lane22_strm1_tmp     ;
  reg [31:0] pe23_lane23_strm0 [0:4095];
  reg [31:0] pe23_lane23_strm0_tmp     ;
  reg [31:0] pe23_lane23_strm1 [0:4095];
  reg [31:0] pe23_lane23_strm1_tmp     ;
  reg [31:0] pe23_lane24_strm0 [0:4095];
  reg [31:0] pe23_lane24_strm0_tmp     ;
  reg [31:0] pe23_lane24_strm1 [0:4095];
  reg [31:0] pe23_lane24_strm1_tmp     ;
  reg [31:0] pe23_lane25_strm0 [0:4095];
  reg [31:0] pe23_lane25_strm0_tmp     ;
  reg [31:0] pe23_lane25_strm1 [0:4095];
  reg [31:0] pe23_lane25_strm1_tmp     ;
  reg [31:0] pe23_lane26_strm0 [0:4095];
  reg [31:0] pe23_lane26_strm0_tmp     ;
  reg [31:0] pe23_lane26_strm1 [0:4095];
  reg [31:0] pe23_lane26_strm1_tmp     ;
  reg [31:0] pe23_lane27_strm0 [0:4095];
  reg [31:0] pe23_lane27_strm0_tmp     ;
  reg [31:0] pe23_lane27_strm1 [0:4095];
  reg [31:0] pe23_lane27_strm1_tmp     ;
  reg [31:0] pe23_lane28_strm0 [0:4095];
  reg [31:0] pe23_lane28_strm0_tmp     ;
  reg [31:0] pe23_lane28_strm1 [0:4095];
  reg [31:0] pe23_lane28_strm1_tmp     ;
  reg [31:0] pe23_lane29_strm0 [0:4095];
  reg [31:0] pe23_lane29_strm0_tmp     ;
  reg [31:0] pe23_lane29_strm1 [0:4095];
  reg [31:0] pe23_lane29_strm1_tmp     ;
  reg [31:0] pe23_lane30_strm0 [0:4095];
  reg [31:0] pe23_lane30_strm0_tmp     ;
  reg [31:0] pe23_lane30_strm1 [0:4095];
  reg [31:0] pe23_lane30_strm1_tmp     ;
  reg [31:0] pe23_lane31_strm0 [0:4095];
  reg [31:0] pe23_lane31_strm0_tmp     ;
  reg [31:0] pe23_lane31_strm1 [0:4095];
  reg [31:0] pe23_lane31_strm1_tmp     ;
  reg [31:0] pe24_lane0_strm0 [0:4095];
  reg [31:0] pe24_lane0_strm0_tmp     ;
  reg [31:0] pe24_lane0_strm1 [0:4095];
  reg [31:0] pe24_lane0_strm1_tmp     ;
  reg [31:0] pe24_lane1_strm0 [0:4095];
  reg [31:0] pe24_lane1_strm0_tmp     ;
  reg [31:0] pe24_lane1_strm1 [0:4095];
  reg [31:0] pe24_lane1_strm1_tmp     ;
  reg [31:0] pe24_lane2_strm0 [0:4095];
  reg [31:0] pe24_lane2_strm0_tmp     ;
  reg [31:0] pe24_lane2_strm1 [0:4095];
  reg [31:0] pe24_lane2_strm1_tmp     ;
  reg [31:0] pe24_lane3_strm0 [0:4095];
  reg [31:0] pe24_lane3_strm0_tmp     ;
  reg [31:0] pe24_lane3_strm1 [0:4095];
  reg [31:0] pe24_lane3_strm1_tmp     ;
  reg [31:0] pe24_lane4_strm0 [0:4095];
  reg [31:0] pe24_lane4_strm0_tmp     ;
  reg [31:0] pe24_lane4_strm1 [0:4095];
  reg [31:0] pe24_lane4_strm1_tmp     ;
  reg [31:0] pe24_lane5_strm0 [0:4095];
  reg [31:0] pe24_lane5_strm0_tmp     ;
  reg [31:0] pe24_lane5_strm1 [0:4095];
  reg [31:0] pe24_lane5_strm1_tmp     ;
  reg [31:0] pe24_lane6_strm0 [0:4095];
  reg [31:0] pe24_lane6_strm0_tmp     ;
  reg [31:0] pe24_lane6_strm1 [0:4095];
  reg [31:0] pe24_lane6_strm1_tmp     ;
  reg [31:0] pe24_lane7_strm0 [0:4095];
  reg [31:0] pe24_lane7_strm0_tmp     ;
  reg [31:0] pe24_lane7_strm1 [0:4095];
  reg [31:0] pe24_lane7_strm1_tmp     ;
  reg [31:0] pe24_lane8_strm0 [0:4095];
  reg [31:0] pe24_lane8_strm0_tmp     ;
  reg [31:0] pe24_lane8_strm1 [0:4095];
  reg [31:0] pe24_lane8_strm1_tmp     ;
  reg [31:0] pe24_lane9_strm0 [0:4095];
  reg [31:0] pe24_lane9_strm0_tmp     ;
  reg [31:0] pe24_lane9_strm1 [0:4095];
  reg [31:0] pe24_lane9_strm1_tmp     ;
  reg [31:0] pe24_lane10_strm0 [0:4095];
  reg [31:0] pe24_lane10_strm0_tmp     ;
  reg [31:0] pe24_lane10_strm1 [0:4095];
  reg [31:0] pe24_lane10_strm1_tmp     ;
  reg [31:0] pe24_lane11_strm0 [0:4095];
  reg [31:0] pe24_lane11_strm0_tmp     ;
  reg [31:0] pe24_lane11_strm1 [0:4095];
  reg [31:0] pe24_lane11_strm1_tmp     ;
  reg [31:0] pe24_lane12_strm0 [0:4095];
  reg [31:0] pe24_lane12_strm0_tmp     ;
  reg [31:0] pe24_lane12_strm1 [0:4095];
  reg [31:0] pe24_lane12_strm1_tmp     ;
  reg [31:0] pe24_lane13_strm0 [0:4095];
  reg [31:0] pe24_lane13_strm0_tmp     ;
  reg [31:0] pe24_lane13_strm1 [0:4095];
  reg [31:0] pe24_lane13_strm1_tmp     ;
  reg [31:0] pe24_lane14_strm0 [0:4095];
  reg [31:0] pe24_lane14_strm0_tmp     ;
  reg [31:0] pe24_lane14_strm1 [0:4095];
  reg [31:0] pe24_lane14_strm1_tmp     ;
  reg [31:0] pe24_lane15_strm0 [0:4095];
  reg [31:0] pe24_lane15_strm0_tmp     ;
  reg [31:0] pe24_lane15_strm1 [0:4095];
  reg [31:0] pe24_lane15_strm1_tmp     ;
  reg [31:0] pe24_lane16_strm0 [0:4095];
  reg [31:0] pe24_lane16_strm0_tmp     ;
  reg [31:0] pe24_lane16_strm1 [0:4095];
  reg [31:0] pe24_lane16_strm1_tmp     ;
  reg [31:0] pe24_lane17_strm0 [0:4095];
  reg [31:0] pe24_lane17_strm0_tmp     ;
  reg [31:0] pe24_lane17_strm1 [0:4095];
  reg [31:0] pe24_lane17_strm1_tmp     ;
  reg [31:0] pe24_lane18_strm0 [0:4095];
  reg [31:0] pe24_lane18_strm0_tmp     ;
  reg [31:0] pe24_lane18_strm1 [0:4095];
  reg [31:0] pe24_lane18_strm1_tmp     ;
  reg [31:0] pe24_lane19_strm0 [0:4095];
  reg [31:0] pe24_lane19_strm0_tmp     ;
  reg [31:0] pe24_lane19_strm1 [0:4095];
  reg [31:0] pe24_lane19_strm1_tmp     ;
  reg [31:0] pe24_lane20_strm0 [0:4095];
  reg [31:0] pe24_lane20_strm0_tmp     ;
  reg [31:0] pe24_lane20_strm1 [0:4095];
  reg [31:0] pe24_lane20_strm1_tmp     ;
  reg [31:0] pe24_lane21_strm0 [0:4095];
  reg [31:0] pe24_lane21_strm0_tmp     ;
  reg [31:0] pe24_lane21_strm1 [0:4095];
  reg [31:0] pe24_lane21_strm1_tmp     ;
  reg [31:0] pe24_lane22_strm0 [0:4095];
  reg [31:0] pe24_lane22_strm0_tmp     ;
  reg [31:0] pe24_lane22_strm1 [0:4095];
  reg [31:0] pe24_lane22_strm1_tmp     ;
  reg [31:0] pe24_lane23_strm0 [0:4095];
  reg [31:0] pe24_lane23_strm0_tmp     ;
  reg [31:0] pe24_lane23_strm1 [0:4095];
  reg [31:0] pe24_lane23_strm1_tmp     ;
  reg [31:0] pe24_lane24_strm0 [0:4095];
  reg [31:0] pe24_lane24_strm0_tmp     ;
  reg [31:0] pe24_lane24_strm1 [0:4095];
  reg [31:0] pe24_lane24_strm1_tmp     ;
  reg [31:0] pe24_lane25_strm0 [0:4095];
  reg [31:0] pe24_lane25_strm0_tmp     ;
  reg [31:0] pe24_lane25_strm1 [0:4095];
  reg [31:0] pe24_lane25_strm1_tmp     ;
  reg [31:0] pe24_lane26_strm0 [0:4095];
  reg [31:0] pe24_lane26_strm0_tmp     ;
  reg [31:0] pe24_lane26_strm1 [0:4095];
  reg [31:0] pe24_lane26_strm1_tmp     ;
  reg [31:0] pe24_lane27_strm0 [0:4095];
  reg [31:0] pe24_lane27_strm0_tmp     ;
  reg [31:0] pe24_lane27_strm1 [0:4095];
  reg [31:0] pe24_lane27_strm1_tmp     ;
  reg [31:0] pe24_lane28_strm0 [0:4095];
  reg [31:0] pe24_lane28_strm0_tmp     ;
  reg [31:0] pe24_lane28_strm1 [0:4095];
  reg [31:0] pe24_lane28_strm1_tmp     ;
  reg [31:0] pe24_lane29_strm0 [0:4095];
  reg [31:0] pe24_lane29_strm0_tmp     ;
  reg [31:0] pe24_lane29_strm1 [0:4095];
  reg [31:0] pe24_lane29_strm1_tmp     ;
  reg [31:0] pe24_lane30_strm0 [0:4095];
  reg [31:0] pe24_lane30_strm0_tmp     ;
  reg [31:0] pe24_lane30_strm1 [0:4095];
  reg [31:0] pe24_lane30_strm1_tmp     ;
  reg [31:0] pe24_lane31_strm0 [0:4095];
  reg [31:0] pe24_lane31_strm0_tmp     ;
  reg [31:0] pe24_lane31_strm1 [0:4095];
  reg [31:0] pe24_lane31_strm1_tmp     ;
  reg [31:0] pe25_lane0_strm0 [0:4095];
  reg [31:0] pe25_lane0_strm0_tmp     ;
  reg [31:0] pe25_lane0_strm1 [0:4095];
  reg [31:0] pe25_lane0_strm1_tmp     ;
  reg [31:0] pe25_lane1_strm0 [0:4095];
  reg [31:0] pe25_lane1_strm0_tmp     ;
  reg [31:0] pe25_lane1_strm1 [0:4095];
  reg [31:0] pe25_lane1_strm1_tmp     ;
  reg [31:0] pe25_lane2_strm0 [0:4095];
  reg [31:0] pe25_lane2_strm0_tmp     ;
  reg [31:0] pe25_lane2_strm1 [0:4095];
  reg [31:0] pe25_lane2_strm1_tmp     ;
  reg [31:0] pe25_lane3_strm0 [0:4095];
  reg [31:0] pe25_lane3_strm0_tmp     ;
  reg [31:0] pe25_lane3_strm1 [0:4095];
  reg [31:0] pe25_lane3_strm1_tmp     ;
  reg [31:0] pe25_lane4_strm0 [0:4095];
  reg [31:0] pe25_lane4_strm0_tmp     ;
  reg [31:0] pe25_lane4_strm1 [0:4095];
  reg [31:0] pe25_lane4_strm1_tmp     ;
  reg [31:0] pe25_lane5_strm0 [0:4095];
  reg [31:0] pe25_lane5_strm0_tmp     ;
  reg [31:0] pe25_lane5_strm1 [0:4095];
  reg [31:0] pe25_lane5_strm1_tmp     ;
  reg [31:0] pe25_lane6_strm0 [0:4095];
  reg [31:0] pe25_lane6_strm0_tmp     ;
  reg [31:0] pe25_lane6_strm1 [0:4095];
  reg [31:0] pe25_lane6_strm1_tmp     ;
  reg [31:0] pe25_lane7_strm0 [0:4095];
  reg [31:0] pe25_lane7_strm0_tmp     ;
  reg [31:0] pe25_lane7_strm1 [0:4095];
  reg [31:0] pe25_lane7_strm1_tmp     ;
  reg [31:0] pe25_lane8_strm0 [0:4095];
  reg [31:0] pe25_lane8_strm0_tmp     ;
  reg [31:0] pe25_lane8_strm1 [0:4095];
  reg [31:0] pe25_lane8_strm1_tmp     ;
  reg [31:0] pe25_lane9_strm0 [0:4095];
  reg [31:0] pe25_lane9_strm0_tmp     ;
  reg [31:0] pe25_lane9_strm1 [0:4095];
  reg [31:0] pe25_lane9_strm1_tmp     ;
  reg [31:0] pe25_lane10_strm0 [0:4095];
  reg [31:0] pe25_lane10_strm0_tmp     ;
  reg [31:0] pe25_lane10_strm1 [0:4095];
  reg [31:0] pe25_lane10_strm1_tmp     ;
  reg [31:0] pe25_lane11_strm0 [0:4095];
  reg [31:0] pe25_lane11_strm0_tmp     ;
  reg [31:0] pe25_lane11_strm1 [0:4095];
  reg [31:0] pe25_lane11_strm1_tmp     ;
  reg [31:0] pe25_lane12_strm0 [0:4095];
  reg [31:0] pe25_lane12_strm0_tmp     ;
  reg [31:0] pe25_lane12_strm1 [0:4095];
  reg [31:0] pe25_lane12_strm1_tmp     ;
  reg [31:0] pe25_lane13_strm0 [0:4095];
  reg [31:0] pe25_lane13_strm0_tmp     ;
  reg [31:0] pe25_lane13_strm1 [0:4095];
  reg [31:0] pe25_lane13_strm1_tmp     ;
  reg [31:0] pe25_lane14_strm0 [0:4095];
  reg [31:0] pe25_lane14_strm0_tmp     ;
  reg [31:0] pe25_lane14_strm1 [0:4095];
  reg [31:0] pe25_lane14_strm1_tmp     ;
  reg [31:0] pe25_lane15_strm0 [0:4095];
  reg [31:0] pe25_lane15_strm0_tmp     ;
  reg [31:0] pe25_lane15_strm1 [0:4095];
  reg [31:0] pe25_lane15_strm1_tmp     ;
  reg [31:0] pe25_lane16_strm0 [0:4095];
  reg [31:0] pe25_lane16_strm0_tmp     ;
  reg [31:0] pe25_lane16_strm1 [0:4095];
  reg [31:0] pe25_lane16_strm1_tmp     ;
  reg [31:0] pe25_lane17_strm0 [0:4095];
  reg [31:0] pe25_lane17_strm0_tmp     ;
  reg [31:0] pe25_lane17_strm1 [0:4095];
  reg [31:0] pe25_lane17_strm1_tmp     ;
  reg [31:0] pe25_lane18_strm0 [0:4095];
  reg [31:0] pe25_lane18_strm0_tmp     ;
  reg [31:0] pe25_lane18_strm1 [0:4095];
  reg [31:0] pe25_lane18_strm1_tmp     ;
  reg [31:0] pe25_lane19_strm0 [0:4095];
  reg [31:0] pe25_lane19_strm0_tmp     ;
  reg [31:0] pe25_lane19_strm1 [0:4095];
  reg [31:0] pe25_lane19_strm1_tmp     ;
  reg [31:0] pe25_lane20_strm0 [0:4095];
  reg [31:0] pe25_lane20_strm0_tmp     ;
  reg [31:0] pe25_lane20_strm1 [0:4095];
  reg [31:0] pe25_lane20_strm1_tmp     ;
  reg [31:0] pe25_lane21_strm0 [0:4095];
  reg [31:0] pe25_lane21_strm0_tmp     ;
  reg [31:0] pe25_lane21_strm1 [0:4095];
  reg [31:0] pe25_lane21_strm1_tmp     ;
  reg [31:0] pe25_lane22_strm0 [0:4095];
  reg [31:0] pe25_lane22_strm0_tmp     ;
  reg [31:0] pe25_lane22_strm1 [0:4095];
  reg [31:0] pe25_lane22_strm1_tmp     ;
  reg [31:0] pe25_lane23_strm0 [0:4095];
  reg [31:0] pe25_lane23_strm0_tmp     ;
  reg [31:0] pe25_lane23_strm1 [0:4095];
  reg [31:0] pe25_lane23_strm1_tmp     ;
  reg [31:0] pe25_lane24_strm0 [0:4095];
  reg [31:0] pe25_lane24_strm0_tmp     ;
  reg [31:0] pe25_lane24_strm1 [0:4095];
  reg [31:0] pe25_lane24_strm1_tmp     ;
  reg [31:0] pe25_lane25_strm0 [0:4095];
  reg [31:0] pe25_lane25_strm0_tmp     ;
  reg [31:0] pe25_lane25_strm1 [0:4095];
  reg [31:0] pe25_lane25_strm1_tmp     ;
  reg [31:0] pe25_lane26_strm0 [0:4095];
  reg [31:0] pe25_lane26_strm0_tmp     ;
  reg [31:0] pe25_lane26_strm1 [0:4095];
  reg [31:0] pe25_lane26_strm1_tmp     ;
  reg [31:0] pe25_lane27_strm0 [0:4095];
  reg [31:0] pe25_lane27_strm0_tmp     ;
  reg [31:0] pe25_lane27_strm1 [0:4095];
  reg [31:0] pe25_lane27_strm1_tmp     ;
  reg [31:0] pe25_lane28_strm0 [0:4095];
  reg [31:0] pe25_lane28_strm0_tmp     ;
  reg [31:0] pe25_lane28_strm1 [0:4095];
  reg [31:0] pe25_lane28_strm1_tmp     ;
  reg [31:0] pe25_lane29_strm0 [0:4095];
  reg [31:0] pe25_lane29_strm0_tmp     ;
  reg [31:0] pe25_lane29_strm1 [0:4095];
  reg [31:0] pe25_lane29_strm1_tmp     ;
  reg [31:0] pe25_lane30_strm0 [0:4095];
  reg [31:0] pe25_lane30_strm0_tmp     ;
  reg [31:0] pe25_lane30_strm1 [0:4095];
  reg [31:0] pe25_lane30_strm1_tmp     ;
  reg [31:0] pe25_lane31_strm0 [0:4095];
  reg [31:0] pe25_lane31_strm0_tmp     ;
  reg [31:0] pe25_lane31_strm1 [0:4095];
  reg [31:0] pe25_lane31_strm1_tmp     ;
  reg [31:0] pe26_lane0_strm0 [0:4095];
  reg [31:0] pe26_lane0_strm0_tmp     ;
  reg [31:0] pe26_lane0_strm1 [0:4095];
  reg [31:0] pe26_lane0_strm1_tmp     ;
  reg [31:0] pe26_lane1_strm0 [0:4095];
  reg [31:0] pe26_lane1_strm0_tmp     ;
  reg [31:0] pe26_lane1_strm1 [0:4095];
  reg [31:0] pe26_lane1_strm1_tmp     ;
  reg [31:0] pe26_lane2_strm0 [0:4095];
  reg [31:0] pe26_lane2_strm0_tmp     ;
  reg [31:0] pe26_lane2_strm1 [0:4095];
  reg [31:0] pe26_lane2_strm1_tmp     ;
  reg [31:0] pe26_lane3_strm0 [0:4095];
  reg [31:0] pe26_lane3_strm0_tmp     ;
  reg [31:0] pe26_lane3_strm1 [0:4095];
  reg [31:0] pe26_lane3_strm1_tmp     ;
  reg [31:0] pe26_lane4_strm0 [0:4095];
  reg [31:0] pe26_lane4_strm0_tmp     ;
  reg [31:0] pe26_lane4_strm1 [0:4095];
  reg [31:0] pe26_lane4_strm1_tmp     ;
  reg [31:0] pe26_lane5_strm0 [0:4095];
  reg [31:0] pe26_lane5_strm0_tmp     ;
  reg [31:0] pe26_lane5_strm1 [0:4095];
  reg [31:0] pe26_lane5_strm1_tmp     ;
  reg [31:0] pe26_lane6_strm0 [0:4095];
  reg [31:0] pe26_lane6_strm0_tmp     ;
  reg [31:0] pe26_lane6_strm1 [0:4095];
  reg [31:0] pe26_lane6_strm1_tmp     ;
  reg [31:0] pe26_lane7_strm0 [0:4095];
  reg [31:0] pe26_lane7_strm0_tmp     ;
  reg [31:0] pe26_lane7_strm1 [0:4095];
  reg [31:0] pe26_lane7_strm1_tmp     ;
  reg [31:0] pe26_lane8_strm0 [0:4095];
  reg [31:0] pe26_lane8_strm0_tmp     ;
  reg [31:0] pe26_lane8_strm1 [0:4095];
  reg [31:0] pe26_lane8_strm1_tmp     ;
  reg [31:0] pe26_lane9_strm0 [0:4095];
  reg [31:0] pe26_lane9_strm0_tmp     ;
  reg [31:0] pe26_lane9_strm1 [0:4095];
  reg [31:0] pe26_lane9_strm1_tmp     ;
  reg [31:0] pe26_lane10_strm0 [0:4095];
  reg [31:0] pe26_lane10_strm0_tmp     ;
  reg [31:0] pe26_lane10_strm1 [0:4095];
  reg [31:0] pe26_lane10_strm1_tmp     ;
  reg [31:0] pe26_lane11_strm0 [0:4095];
  reg [31:0] pe26_lane11_strm0_tmp     ;
  reg [31:0] pe26_lane11_strm1 [0:4095];
  reg [31:0] pe26_lane11_strm1_tmp     ;
  reg [31:0] pe26_lane12_strm0 [0:4095];
  reg [31:0] pe26_lane12_strm0_tmp     ;
  reg [31:0] pe26_lane12_strm1 [0:4095];
  reg [31:0] pe26_lane12_strm1_tmp     ;
  reg [31:0] pe26_lane13_strm0 [0:4095];
  reg [31:0] pe26_lane13_strm0_tmp     ;
  reg [31:0] pe26_lane13_strm1 [0:4095];
  reg [31:0] pe26_lane13_strm1_tmp     ;
  reg [31:0] pe26_lane14_strm0 [0:4095];
  reg [31:0] pe26_lane14_strm0_tmp     ;
  reg [31:0] pe26_lane14_strm1 [0:4095];
  reg [31:0] pe26_lane14_strm1_tmp     ;
  reg [31:0] pe26_lane15_strm0 [0:4095];
  reg [31:0] pe26_lane15_strm0_tmp     ;
  reg [31:0] pe26_lane15_strm1 [0:4095];
  reg [31:0] pe26_lane15_strm1_tmp     ;
  reg [31:0] pe26_lane16_strm0 [0:4095];
  reg [31:0] pe26_lane16_strm0_tmp     ;
  reg [31:0] pe26_lane16_strm1 [0:4095];
  reg [31:0] pe26_lane16_strm1_tmp     ;
  reg [31:0] pe26_lane17_strm0 [0:4095];
  reg [31:0] pe26_lane17_strm0_tmp     ;
  reg [31:0] pe26_lane17_strm1 [0:4095];
  reg [31:0] pe26_lane17_strm1_tmp     ;
  reg [31:0] pe26_lane18_strm0 [0:4095];
  reg [31:0] pe26_lane18_strm0_tmp     ;
  reg [31:0] pe26_lane18_strm1 [0:4095];
  reg [31:0] pe26_lane18_strm1_tmp     ;
  reg [31:0] pe26_lane19_strm0 [0:4095];
  reg [31:0] pe26_lane19_strm0_tmp     ;
  reg [31:0] pe26_lane19_strm1 [0:4095];
  reg [31:0] pe26_lane19_strm1_tmp     ;
  reg [31:0] pe26_lane20_strm0 [0:4095];
  reg [31:0] pe26_lane20_strm0_tmp     ;
  reg [31:0] pe26_lane20_strm1 [0:4095];
  reg [31:0] pe26_lane20_strm1_tmp     ;
  reg [31:0] pe26_lane21_strm0 [0:4095];
  reg [31:0] pe26_lane21_strm0_tmp     ;
  reg [31:0] pe26_lane21_strm1 [0:4095];
  reg [31:0] pe26_lane21_strm1_tmp     ;
  reg [31:0] pe26_lane22_strm0 [0:4095];
  reg [31:0] pe26_lane22_strm0_tmp     ;
  reg [31:0] pe26_lane22_strm1 [0:4095];
  reg [31:0] pe26_lane22_strm1_tmp     ;
  reg [31:0] pe26_lane23_strm0 [0:4095];
  reg [31:0] pe26_lane23_strm0_tmp     ;
  reg [31:0] pe26_lane23_strm1 [0:4095];
  reg [31:0] pe26_lane23_strm1_tmp     ;
  reg [31:0] pe26_lane24_strm0 [0:4095];
  reg [31:0] pe26_lane24_strm0_tmp     ;
  reg [31:0] pe26_lane24_strm1 [0:4095];
  reg [31:0] pe26_lane24_strm1_tmp     ;
  reg [31:0] pe26_lane25_strm0 [0:4095];
  reg [31:0] pe26_lane25_strm0_tmp     ;
  reg [31:0] pe26_lane25_strm1 [0:4095];
  reg [31:0] pe26_lane25_strm1_tmp     ;
  reg [31:0] pe26_lane26_strm0 [0:4095];
  reg [31:0] pe26_lane26_strm0_tmp     ;
  reg [31:0] pe26_lane26_strm1 [0:4095];
  reg [31:0] pe26_lane26_strm1_tmp     ;
  reg [31:0] pe26_lane27_strm0 [0:4095];
  reg [31:0] pe26_lane27_strm0_tmp     ;
  reg [31:0] pe26_lane27_strm1 [0:4095];
  reg [31:0] pe26_lane27_strm1_tmp     ;
  reg [31:0] pe26_lane28_strm0 [0:4095];
  reg [31:0] pe26_lane28_strm0_tmp     ;
  reg [31:0] pe26_lane28_strm1 [0:4095];
  reg [31:0] pe26_lane28_strm1_tmp     ;
  reg [31:0] pe26_lane29_strm0 [0:4095];
  reg [31:0] pe26_lane29_strm0_tmp     ;
  reg [31:0] pe26_lane29_strm1 [0:4095];
  reg [31:0] pe26_lane29_strm1_tmp     ;
  reg [31:0] pe26_lane30_strm0 [0:4095];
  reg [31:0] pe26_lane30_strm0_tmp     ;
  reg [31:0] pe26_lane30_strm1 [0:4095];
  reg [31:0] pe26_lane30_strm1_tmp     ;
  reg [31:0] pe26_lane31_strm0 [0:4095];
  reg [31:0] pe26_lane31_strm0_tmp     ;
  reg [31:0] pe26_lane31_strm1 [0:4095];
  reg [31:0] pe26_lane31_strm1_tmp     ;
  reg [31:0] pe27_lane0_strm0 [0:4095];
  reg [31:0] pe27_lane0_strm0_tmp     ;
  reg [31:0] pe27_lane0_strm1 [0:4095];
  reg [31:0] pe27_lane0_strm1_tmp     ;
  reg [31:0] pe27_lane1_strm0 [0:4095];
  reg [31:0] pe27_lane1_strm0_tmp     ;
  reg [31:0] pe27_lane1_strm1 [0:4095];
  reg [31:0] pe27_lane1_strm1_tmp     ;
  reg [31:0] pe27_lane2_strm0 [0:4095];
  reg [31:0] pe27_lane2_strm0_tmp     ;
  reg [31:0] pe27_lane2_strm1 [0:4095];
  reg [31:0] pe27_lane2_strm1_tmp     ;
  reg [31:0] pe27_lane3_strm0 [0:4095];
  reg [31:0] pe27_lane3_strm0_tmp     ;
  reg [31:0] pe27_lane3_strm1 [0:4095];
  reg [31:0] pe27_lane3_strm1_tmp     ;
  reg [31:0] pe27_lane4_strm0 [0:4095];
  reg [31:0] pe27_lane4_strm0_tmp     ;
  reg [31:0] pe27_lane4_strm1 [0:4095];
  reg [31:0] pe27_lane4_strm1_tmp     ;
  reg [31:0] pe27_lane5_strm0 [0:4095];
  reg [31:0] pe27_lane5_strm0_tmp     ;
  reg [31:0] pe27_lane5_strm1 [0:4095];
  reg [31:0] pe27_lane5_strm1_tmp     ;
  reg [31:0] pe27_lane6_strm0 [0:4095];
  reg [31:0] pe27_lane6_strm0_tmp     ;
  reg [31:0] pe27_lane6_strm1 [0:4095];
  reg [31:0] pe27_lane6_strm1_tmp     ;
  reg [31:0] pe27_lane7_strm0 [0:4095];
  reg [31:0] pe27_lane7_strm0_tmp     ;
  reg [31:0] pe27_lane7_strm1 [0:4095];
  reg [31:0] pe27_lane7_strm1_tmp     ;
  reg [31:0] pe27_lane8_strm0 [0:4095];
  reg [31:0] pe27_lane8_strm0_tmp     ;
  reg [31:0] pe27_lane8_strm1 [0:4095];
  reg [31:0] pe27_lane8_strm1_tmp     ;
  reg [31:0] pe27_lane9_strm0 [0:4095];
  reg [31:0] pe27_lane9_strm0_tmp     ;
  reg [31:0] pe27_lane9_strm1 [0:4095];
  reg [31:0] pe27_lane9_strm1_tmp     ;
  reg [31:0] pe27_lane10_strm0 [0:4095];
  reg [31:0] pe27_lane10_strm0_tmp     ;
  reg [31:0] pe27_lane10_strm1 [0:4095];
  reg [31:0] pe27_lane10_strm1_tmp     ;
  reg [31:0] pe27_lane11_strm0 [0:4095];
  reg [31:0] pe27_lane11_strm0_tmp     ;
  reg [31:0] pe27_lane11_strm1 [0:4095];
  reg [31:0] pe27_lane11_strm1_tmp     ;
  reg [31:0] pe27_lane12_strm0 [0:4095];
  reg [31:0] pe27_lane12_strm0_tmp     ;
  reg [31:0] pe27_lane12_strm1 [0:4095];
  reg [31:0] pe27_lane12_strm1_tmp     ;
  reg [31:0] pe27_lane13_strm0 [0:4095];
  reg [31:0] pe27_lane13_strm0_tmp     ;
  reg [31:0] pe27_lane13_strm1 [0:4095];
  reg [31:0] pe27_lane13_strm1_tmp     ;
  reg [31:0] pe27_lane14_strm0 [0:4095];
  reg [31:0] pe27_lane14_strm0_tmp     ;
  reg [31:0] pe27_lane14_strm1 [0:4095];
  reg [31:0] pe27_lane14_strm1_tmp     ;
  reg [31:0] pe27_lane15_strm0 [0:4095];
  reg [31:0] pe27_lane15_strm0_tmp     ;
  reg [31:0] pe27_lane15_strm1 [0:4095];
  reg [31:0] pe27_lane15_strm1_tmp     ;
  reg [31:0] pe27_lane16_strm0 [0:4095];
  reg [31:0] pe27_lane16_strm0_tmp     ;
  reg [31:0] pe27_lane16_strm1 [0:4095];
  reg [31:0] pe27_lane16_strm1_tmp     ;
  reg [31:0] pe27_lane17_strm0 [0:4095];
  reg [31:0] pe27_lane17_strm0_tmp     ;
  reg [31:0] pe27_lane17_strm1 [0:4095];
  reg [31:0] pe27_lane17_strm1_tmp     ;
  reg [31:0] pe27_lane18_strm0 [0:4095];
  reg [31:0] pe27_lane18_strm0_tmp     ;
  reg [31:0] pe27_lane18_strm1 [0:4095];
  reg [31:0] pe27_lane18_strm1_tmp     ;
  reg [31:0] pe27_lane19_strm0 [0:4095];
  reg [31:0] pe27_lane19_strm0_tmp     ;
  reg [31:0] pe27_lane19_strm1 [0:4095];
  reg [31:0] pe27_lane19_strm1_tmp     ;
  reg [31:0] pe27_lane20_strm0 [0:4095];
  reg [31:0] pe27_lane20_strm0_tmp     ;
  reg [31:0] pe27_lane20_strm1 [0:4095];
  reg [31:0] pe27_lane20_strm1_tmp     ;
  reg [31:0] pe27_lane21_strm0 [0:4095];
  reg [31:0] pe27_lane21_strm0_tmp     ;
  reg [31:0] pe27_lane21_strm1 [0:4095];
  reg [31:0] pe27_lane21_strm1_tmp     ;
  reg [31:0] pe27_lane22_strm0 [0:4095];
  reg [31:0] pe27_lane22_strm0_tmp     ;
  reg [31:0] pe27_lane22_strm1 [0:4095];
  reg [31:0] pe27_lane22_strm1_tmp     ;
  reg [31:0] pe27_lane23_strm0 [0:4095];
  reg [31:0] pe27_lane23_strm0_tmp     ;
  reg [31:0] pe27_lane23_strm1 [0:4095];
  reg [31:0] pe27_lane23_strm1_tmp     ;
  reg [31:0] pe27_lane24_strm0 [0:4095];
  reg [31:0] pe27_lane24_strm0_tmp     ;
  reg [31:0] pe27_lane24_strm1 [0:4095];
  reg [31:0] pe27_lane24_strm1_tmp     ;
  reg [31:0] pe27_lane25_strm0 [0:4095];
  reg [31:0] pe27_lane25_strm0_tmp     ;
  reg [31:0] pe27_lane25_strm1 [0:4095];
  reg [31:0] pe27_lane25_strm1_tmp     ;
  reg [31:0] pe27_lane26_strm0 [0:4095];
  reg [31:0] pe27_lane26_strm0_tmp     ;
  reg [31:0] pe27_lane26_strm1 [0:4095];
  reg [31:0] pe27_lane26_strm1_tmp     ;
  reg [31:0] pe27_lane27_strm0 [0:4095];
  reg [31:0] pe27_lane27_strm0_tmp     ;
  reg [31:0] pe27_lane27_strm1 [0:4095];
  reg [31:0] pe27_lane27_strm1_tmp     ;
  reg [31:0] pe27_lane28_strm0 [0:4095];
  reg [31:0] pe27_lane28_strm0_tmp     ;
  reg [31:0] pe27_lane28_strm1 [0:4095];
  reg [31:0] pe27_lane28_strm1_tmp     ;
  reg [31:0] pe27_lane29_strm0 [0:4095];
  reg [31:0] pe27_lane29_strm0_tmp     ;
  reg [31:0] pe27_lane29_strm1 [0:4095];
  reg [31:0] pe27_lane29_strm1_tmp     ;
  reg [31:0] pe27_lane30_strm0 [0:4095];
  reg [31:0] pe27_lane30_strm0_tmp     ;
  reg [31:0] pe27_lane30_strm1 [0:4095];
  reg [31:0] pe27_lane30_strm1_tmp     ;
  reg [31:0] pe27_lane31_strm0 [0:4095];
  reg [31:0] pe27_lane31_strm0_tmp     ;
  reg [31:0] pe27_lane31_strm1 [0:4095];
  reg [31:0] pe27_lane31_strm1_tmp     ;
  reg [31:0] pe28_lane0_strm0 [0:4095];
  reg [31:0] pe28_lane0_strm0_tmp     ;
  reg [31:0] pe28_lane0_strm1 [0:4095];
  reg [31:0] pe28_lane0_strm1_tmp     ;
  reg [31:0] pe28_lane1_strm0 [0:4095];
  reg [31:0] pe28_lane1_strm0_tmp     ;
  reg [31:0] pe28_lane1_strm1 [0:4095];
  reg [31:0] pe28_lane1_strm1_tmp     ;
  reg [31:0] pe28_lane2_strm0 [0:4095];
  reg [31:0] pe28_lane2_strm0_tmp     ;
  reg [31:0] pe28_lane2_strm1 [0:4095];
  reg [31:0] pe28_lane2_strm1_tmp     ;
  reg [31:0] pe28_lane3_strm0 [0:4095];
  reg [31:0] pe28_lane3_strm0_tmp     ;
  reg [31:0] pe28_lane3_strm1 [0:4095];
  reg [31:0] pe28_lane3_strm1_tmp     ;
  reg [31:0] pe28_lane4_strm0 [0:4095];
  reg [31:0] pe28_lane4_strm0_tmp     ;
  reg [31:0] pe28_lane4_strm1 [0:4095];
  reg [31:0] pe28_lane4_strm1_tmp     ;
  reg [31:0] pe28_lane5_strm0 [0:4095];
  reg [31:0] pe28_lane5_strm0_tmp     ;
  reg [31:0] pe28_lane5_strm1 [0:4095];
  reg [31:0] pe28_lane5_strm1_tmp     ;
  reg [31:0] pe28_lane6_strm0 [0:4095];
  reg [31:0] pe28_lane6_strm0_tmp     ;
  reg [31:0] pe28_lane6_strm1 [0:4095];
  reg [31:0] pe28_lane6_strm1_tmp     ;
  reg [31:0] pe28_lane7_strm0 [0:4095];
  reg [31:0] pe28_lane7_strm0_tmp     ;
  reg [31:0] pe28_lane7_strm1 [0:4095];
  reg [31:0] pe28_lane7_strm1_tmp     ;
  reg [31:0] pe28_lane8_strm0 [0:4095];
  reg [31:0] pe28_lane8_strm0_tmp     ;
  reg [31:0] pe28_lane8_strm1 [0:4095];
  reg [31:0] pe28_lane8_strm1_tmp     ;
  reg [31:0] pe28_lane9_strm0 [0:4095];
  reg [31:0] pe28_lane9_strm0_tmp     ;
  reg [31:0] pe28_lane9_strm1 [0:4095];
  reg [31:0] pe28_lane9_strm1_tmp     ;
  reg [31:0] pe28_lane10_strm0 [0:4095];
  reg [31:0] pe28_lane10_strm0_tmp     ;
  reg [31:0] pe28_lane10_strm1 [0:4095];
  reg [31:0] pe28_lane10_strm1_tmp     ;
  reg [31:0] pe28_lane11_strm0 [0:4095];
  reg [31:0] pe28_lane11_strm0_tmp     ;
  reg [31:0] pe28_lane11_strm1 [0:4095];
  reg [31:0] pe28_lane11_strm1_tmp     ;
  reg [31:0] pe28_lane12_strm0 [0:4095];
  reg [31:0] pe28_lane12_strm0_tmp     ;
  reg [31:0] pe28_lane12_strm1 [0:4095];
  reg [31:0] pe28_lane12_strm1_tmp     ;
  reg [31:0] pe28_lane13_strm0 [0:4095];
  reg [31:0] pe28_lane13_strm0_tmp     ;
  reg [31:0] pe28_lane13_strm1 [0:4095];
  reg [31:0] pe28_lane13_strm1_tmp     ;
  reg [31:0] pe28_lane14_strm0 [0:4095];
  reg [31:0] pe28_lane14_strm0_tmp     ;
  reg [31:0] pe28_lane14_strm1 [0:4095];
  reg [31:0] pe28_lane14_strm1_tmp     ;
  reg [31:0] pe28_lane15_strm0 [0:4095];
  reg [31:0] pe28_lane15_strm0_tmp     ;
  reg [31:0] pe28_lane15_strm1 [0:4095];
  reg [31:0] pe28_lane15_strm1_tmp     ;
  reg [31:0] pe28_lane16_strm0 [0:4095];
  reg [31:0] pe28_lane16_strm0_tmp     ;
  reg [31:0] pe28_lane16_strm1 [0:4095];
  reg [31:0] pe28_lane16_strm1_tmp     ;
  reg [31:0] pe28_lane17_strm0 [0:4095];
  reg [31:0] pe28_lane17_strm0_tmp     ;
  reg [31:0] pe28_lane17_strm1 [0:4095];
  reg [31:0] pe28_lane17_strm1_tmp     ;
  reg [31:0] pe28_lane18_strm0 [0:4095];
  reg [31:0] pe28_lane18_strm0_tmp     ;
  reg [31:0] pe28_lane18_strm1 [0:4095];
  reg [31:0] pe28_lane18_strm1_tmp     ;
  reg [31:0] pe28_lane19_strm0 [0:4095];
  reg [31:0] pe28_lane19_strm0_tmp     ;
  reg [31:0] pe28_lane19_strm1 [0:4095];
  reg [31:0] pe28_lane19_strm1_tmp     ;
  reg [31:0] pe28_lane20_strm0 [0:4095];
  reg [31:0] pe28_lane20_strm0_tmp     ;
  reg [31:0] pe28_lane20_strm1 [0:4095];
  reg [31:0] pe28_lane20_strm1_tmp     ;
  reg [31:0] pe28_lane21_strm0 [0:4095];
  reg [31:0] pe28_lane21_strm0_tmp     ;
  reg [31:0] pe28_lane21_strm1 [0:4095];
  reg [31:0] pe28_lane21_strm1_tmp     ;
  reg [31:0] pe28_lane22_strm0 [0:4095];
  reg [31:0] pe28_lane22_strm0_tmp     ;
  reg [31:0] pe28_lane22_strm1 [0:4095];
  reg [31:0] pe28_lane22_strm1_tmp     ;
  reg [31:0] pe28_lane23_strm0 [0:4095];
  reg [31:0] pe28_lane23_strm0_tmp     ;
  reg [31:0] pe28_lane23_strm1 [0:4095];
  reg [31:0] pe28_lane23_strm1_tmp     ;
  reg [31:0] pe28_lane24_strm0 [0:4095];
  reg [31:0] pe28_lane24_strm0_tmp     ;
  reg [31:0] pe28_lane24_strm1 [0:4095];
  reg [31:0] pe28_lane24_strm1_tmp     ;
  reg [31:0] pe28_lane25_strm0 [0:4095];
  reg [31:0] pe28_lane25_strm0_tmp     ;
  reg [31:0] pe28_lane25_strm1 [0:4095];
  reg [31:0] pe28_lane25_strm1_tmp     ;
  reg [31:0] pe28_lane26_strm0 [0:4095];
  reg [31:0] pe28_lane26_strm0_tmp     ;
  reg [31:0] pe28_lane26_strm1 [0:4095];
  reg [31:0] pe28_lane26_strm1_tmp     ;
  reg [31:0] pe28_lane27_strm0 [0:4095];
  reg [31:0] pe28_lane27_strm0_tmp     ;
  reg [31:0] pe28_lane27_strm1 [0:4095];
  reg [31:0] pe28_lane27_strm1_tmp     ;
  reg [31:0] pe28_lane28_strm0 [0:4095];
  reg [31:0] pe28_lane28_strm0_tmp     ;
  reg [31:0] pe28_lane28_strm1 [0:4095];
  reg [31:0] pe28_lane28_strm1_tmp     ;
  reg [31:0] pe28_lane29_strm0 [0:4095];
  reg [31:0] pe28_lane29_strm0_tmp     ;
  reg [31:0] pe28_lane29_strm1 [0:4095];
  reg [31:0] pe28_lane29_strm1_tmp     ;
  reg [31:0] pe28_lane30_strm0 [0:4095];
  reg [31:0] pe28_lane30_strm0_tmp     ;
  reg [31:0] pe28_lane30_strm1 [0:4095];
  reg [31:0] pe28_lane30_strm1_tmp     ;
  reg [31:0] pe28_lane31_strm0 [0:4095];
  reg [31:0] pe28_lane31_strm0_tmp     ;
  reg [31:0] pe28_lane31_strm1 [0:4095];
  reg [31:0] pe28_lane31_strm1_tmp     ;
  reg [31:0] pe29_lane0_strm0 [0:4095];
  reg [31:0] pe29_lane0_strm0_tmp     ;
  reg [31:0] pe29_lane0_strm1 [0:4095];
  reg [31:0] pe29_lane0_strm1_tmp     ;
  reg [31:0] pe29_lane1_strm0 [0:4095];
  reg [31:0] pe29_lane1_strm0_tmp     ;
  reg [31:0] pe29_lane1_strm1 [0:4095];
  reg [31:0] pe29_lane1_strm1_tmp     ;
  reg [31:0] pe29_lane2_strm0 [0:4095];
  reg [31:0] pe29_lane2_strm0_tmp     ;
  reg [31:0] pe29_lane2_strm1 [0:4095];
  reg [31:0] pe29_lane2_strm1_tmp     ;
  reg [31:0] pe29_lane3_strm0 [0:4095];
  reg [31:0] pe29_lane3_strm0_tmp     ;
  reg [31:0] pe29_lane3_strm1 [0:4095];
  reg [31:0] pe29_lane3_strm1_tmp     ;
  reg [31:0] pe29_lane4_strm0 [0:4095];
  reg [31:0] pe29_lane4_strm0_tmp     ;
  reg [31:0] pe29_lane4_strm1 [0:4095];
  reg [31:0] pe29_lane4_strm1_tmp     ;
  reg [31:0] pe29_lane5_strm0 [0:4095];
  reg [31:0] pe29_lane5_strm0_tmp     ;
  reg [31:0] pe29_lane5_strm1 [0:4095];
  reg [31:0] pe29_lane5_strm1_tmp     ;
  reg [31:0] pe29_lane6_strm0 [0:4095];
  reg [31:0] pe29_lane6_strm0_tmp     ;
  reg [31:0] pe29_lane6_strm1 [0:4095];
  reg [31:0] pe29_lane6_strm1_tmp     ;
  reg [31:0] pe29_lane7_strm0 [0:4095];
  reg [31:0] pe29_lane7_strm0_tmp     ;
  reg [31:0] pe29_lane7_strm1 [0:4095];
  reg [31:0] pe29_lane7_strm1_tmp     ;
  reg [31:0] pe29_lane8_strm0 [0:4095];
  reg [31:0] pe29_lane8_strm0_tmp     ;
  reg [31:0] pe29_lane8_strm1 [0:4095];
  reg [31:0] pe29_lane8_strm1_tmp     ;
  reg [31:0] pe29_lane9_strm0 [0:4095];
  reg [31:0] pe29_lane9_strm0_tmp     ;
  reg [31:0] pe29_lane9_strm1 [0:4095];
  reg [31:0] pe29_lane9_strm1_tmp     ;
  reg [31:0] pe29_lane10_strm0 [0:4095];
  reg [31:0] pe29_lane10_strm0_tmp     ;
  reg [31:0] pe29_lane10_strm1 [0:4095];
  reg [31:0] pe29_lane10_strm1_tmp     ;
  reg [31:0] pe29_lane11_strm0 [0:4095];
  reg [31:0] pe29_lane11_strm0_tmp     ;
  reg [31:0] pe29_lane11_strm1 [0:4095];
  reg [31:0] pe29_lane11_strm1_tmp     ;
  reg [31:0] pe29_lane12_strm0 [0:4095];
  reg [31:0] pe29_lane12_strm0_tmp     ;
  reg [31:0] pe29_lane12_strm1 [0:4095];
  reg [31:0] pe29_lane12_strm1_tmp     ;
  reg [31:0] pe29_lane13_strm0 [0:4095];
  reg [31:0] pe29_lane13_strm0_tmp     ;
  reg [31:0] pe29_lane13_strm1 [0:4095];
  reg [31:0] pe29_lane13_strm1_tmp     ;
  reg [31:0] pe29_lane14_strm0 [0:4095];
  reg [31:0] pe29_lane14_strm0_tmp     ;
  reg [31:0] pe29_lane14_strm1 [0:4095];
  reg [31:0] pe29_lane14_strm1_tmp     ;
  reg [31:0] pe29_lane15_strm0 [0:4095];
  reg [31:0] pe29_lane15_strm0_tmp     ;
  reg [31:0] pe29_lane15_strm1 [0:4095];
  reg [31:0] pe29_lane15_strm1_tmp     ;
  reg [31:0] pe29_lane16_strm0 [0:4095];
  reg [31:0] pe29_lane16_strm0_tmp     ;
  reg [31:0] pe29_lane16_strm1 [0:4095];
  reg [31:0] pe29_lane16_strm1_tmp     ;
  reg [31:0] pe29_lane17_strm0 [0:4095];
  reg [31:0] pe29_lane17_strm0_tmp     ;
  reg [31:0] pe29_lane17_strm1 [0:4095];
  reg [31:0] pe29_lane17_strm1_tmp     ;
  reg [31:0] pe29_lane18_strm0 [0:4095];
  reg [31:0] pe29_lane18_strm0_tmp     ;
  reg [31:0] pe29_lane18_strm1 [0:4095];
  reg [31:0] pe29_lane18_strm1_tmp     ;
  reg [31:0] pe29_lane19_strm0 [0:4095];
  reg [31:0] pe29_lane19_strm0_tmp     ;
  reg [31:0] pe29_lane19_strm1 [0:4095];
  reg [31:0] pe29_lane19_strm1_tmp     ;
  reg [31:0] pe29_lane20_strm0 [0:4095];
  reg [31:0] pe29_lane20_strm0_tmp     ;
  reg [31:0] pe29_lane20_strm1 [0:4095];
  reg [31:0] pe29_lane20_strm1_tmp     ;
  reg [31:0] pe29_lane21_strm0 [0:4095];
  reg [31:0] pe29_lane21_strm0_tmp     ;
  reg [31:0] pe29_lane21_strm1 [0:4095];
  reg [31:0] pe29_lane21_strm1_tmp     ;
  reg [31:0] pe29_lane22_strm0 [0:4095];
  reg [31:0] pe29_lane22_strm0_tmp     ;
  reg [31:0] pe29_lane22_strm1 [0:4095];
  reg [31:0] pe29_lane22_strm1_tmp     ;
  reg [31:0] pe29_lane23_strm0 [0:4095];
  reg [31:0] pe29_lane23_strm0_tmp     ;
  reg [31:0] pe29_lane23_strm1 [0:4095];
  reg [31:0] pe29_lane23_strm1_tmp     ;
  reg [31:0] pe29_lane24_strm0 [0:4095];
  reg [31:0] pe29_lane24_strm0_tmp     ;
  reg [31:0] pe29_lane24_strm1 [0:4095];
  reg [31:0] pe29_lane24_strm1_tmp     ;
  reg [31:0] pe29_lane25_strm0 [0:4095];
  reg [31:0] pe29_lane25_strm0_tmp     ;
  reg [31:0] pe29_lane25_strm1 [0:4095];
  reg [31:0] pe29_lane25_strm1_tmp     ;
  reg [31:0] pe29_lane26_strm0 [0:4095];
  reg [31:0] pe29_lane26_strm0_tmp     ;
  reg [31:0] pe29_lane26_strm1 [0:4095];
  reg [31:0] pe29_lane26_strm1_tmp     ;
  reg [31:0] pe29_lane27_strm0 [0:4095];
  reg [31:0] pe29_lane27_strm0_tmp     ;
  reg [31:0] pe29_lane27_strm1 [0:4095];
  reg [31:0] pe29_lane27_strm1_tmp     ;
  reg [31:0] pe29_lane28_strm0 [0:4095];
  reg [31:0] pe29_lane28_strm0_tmp     ;
  reg [31:0] pe29_lane28_strm1 [0:4095];
  reg [31:0] pe29_lane28_strm1_tmp     ;
  reg [31:0] pe29_lane29_strm0 [0:4095];
  reg [31:0] pe29_lane29_strm0_tmp     ;
  reg [31:0] pe29_lane29_strm1 [0:4095];
  reg [31:0] pe29_lane29_strm1_tmp     ;
  reg [31:0] pe29_lane30_strm0 [0:4095];
  reg [31:0] pe29_lane30_strm0_tmp     ;
  reg [31:0] pe29_lane30_strm1 [0:4095];
  reg [31:0] pe29_lane30_strm1_tmp     ;
  reg [31:0] pe29_lane31_strm0 [0:4095];
  reg [31:0] pe29_lane31_strm0_tmp     ;
  reg [31:0] pe29_lane31_strm1 [0:4095];
  reg [31:0] pe29_lane31_strm1_tmp     ;
  reg [31:0] pe30_lane0_strm0 [0:4095];
  reg [31:0] pe30_lane0_strm0_tmp     ;
  reg [31:0] pe30_lane0_strm1 [0:4095];
  reg [31:0] pe30_lane0_strm1_tmp     ;
  reg [31:0] pe30_lane1_strm0 [0:4095];
  reg [31:0] pe30_lane1_strm0_tmp     ;
  reg [31:0] pe30_lane1_strm1 [0:4095];
  reg [31:0] pe30_lane1_strm1_tmp     ;
  reg [31:0] pe30_lane2_strm0 [0:4095];
  reg [31:0] pe30_lane2_strm0_tmp     ;
  reg [31:0] pe30_lane2_strm1 [0:4095];
  reg [31:0] pe30_lane2_strm1_tmp     ;
  reg [31:0] pe30_lane3_strm0 [0:4095];
  reg [31:0] pe30_lane3_strm0_tmp     ;
  reg [31:0] pe30_lane3_strm1 [0:4095];
  reg [31:0] pe30_lane3_strm1_tmp     ;
  reg [31:0] pe30_lane4_strm0 [0:4095];
  reg [31:0] pe30_lane4_strm0_tmp     ;
  reg [31:0] pe30_lane4_strm1 [0:4095];
  reg [31:0] pe30_lane4_strm1_tmp     ;
  reg [31:0] pe30_lane5_strm0 [0:4095];
  reg [31:0] pe30_lane5_strm0_tmp     ;
  reg [31:0] pe30_lane5_strm1 [0:4095];
  reg [31:0] pe30_lane5_strm1_tmp     ;
  reg [31:0] pe30_lane6_strm0 [0:4095];
  reg [31:0] pe30_lane6_strm0_tmp     ;
  reg [31:0] pe30_lane6_strm1 [0:4095];
  reg [31:0] pe30_lane6_strm1_tmp     ;
  reg [31:0] pe30_lane7_strm0 [0:4095];
  reg [31:0] pe30_lane7_strm0_tmp     ;
  reg [31:0] pe30_lane7_strm1 [0:4095];
  reg [31:0] pe30_lane7_strm1_tmp     ;
  reg [31:0] pe30_lane8_strm0 [0:4095];
  reg [31:0] pe30_lane8_strm0_tmp     ;
  reg [31:0] pe30_lane8_strm1 [0:4095];
  reg [31:0] pe30_lane8_strm1_tmp     ;
  reg [31:0] pe30_lane9_strm0 [0:4095];
  reg [31:0] pe30_lane9_strm0_tmp     ;
  reg [31:0] pe30_lane9_strm1 [0:4095];
  reg [31:0] pe30_lane9_strm1_tmp     ;
  reg [31:0] pe30_lane10_strm0 [0:4095];
  reg [31:0] pe30_lane10_strm0_tmp     ;
  reg [31:0] pe30_lane10_strm1 [0:4095];
  reg [31:0] pe30_lane10_strm1_tmp     ;
  reg [31:0] pe30_lane11_strm0 [0:4095];
  reg [31:0] pe30_lane11_strm0_tmp     ;
  reg [31:0] pe30_lane11_strm1 [0:4095];
  reg [31:0] pe30_lane11_strm1_tmp     ;
  reg [31:0] pe30_lane12_strm0 [0:4095];
  reg [31:0] pe30_lane12_strm0_tmp     ;
  reg [31:0] pe30_lane12_strm1 [0:4095];
  reg [31:0] pe30_lane12_strm1_tmp     ;
  reg [31:0] pe30_lane13_strm0 [0:4095];
  reg [31:0] pe30_lane13_strm0_tmp     ;
  reg [31:0] pe30_lane13_strm1 [0:4095];
  reg [31:0] pe30_lane13_strm1_tmp     ;
  reg [31:0] pe30_lane14_strm0 [0:4095];
  reg [31:0] pe30_lane14_strm0_tmp     ;
  reg [31:0] pe30_lane14_strm1 [0:4095];
  reg [31:0] pe30_lane14_strm1_tmp     ;
  reg [31:0] pe30_lane15_strm0 [0:4095];
  reg [31:0] pe30_lane15_strm0_tmp     ;
  reg [31:0] pe30_lane15_strm1 [0:4095];
  reg [31:0] pe30_lane15_strm1_tmp     ;
  reg [31:0] pe30_lane16_strm0 [0:4095];
  reg [31:0] pe30_lane16_strm0_tmp     ;
  reg [31:0] pe30_lane16_strm1 [0:4095];
  reg [31:0] pe30_lane16_strm1_tmp     ;
  reg [31:0] pe30_lane17_strm0 [0:4095];
  reg [31:0] pe30_lane17_strm0_tmp     ;
  reg [31:0] pe30_lane17_strm1 [0:4095];
  reg [31:0] pe30_lane17_strm1_tmp     ;
  reg [31:0] pe30_lane18_strm0 [0:4095];
  reg [31:0] pe30_lane18_strm0_tmp     ;
  reg [31:0] pe30_lane18_strm1 [0:4095];
  reg [31:0] pe30_lane18_strm1_tmp     ;
  reg [31:0] pe30_lane19_strm0 [0:4095];
  reg [31:0] pe30_lane19_strm0_tmp     ;
  reg [31:0] pe30_lane19_strm1 [0:4095];
  reg [31:0] pe30_lane19_strm1_tmp     ;
  reg [31:0] pe30_lane20_strm0 [0:4095];
  reg [31:0] pe30_lane20_strm0_tmp     ;
  reg [31:0] pe30_lane20_strm1 [0:4095];
  reg [31:0] pe30_lane20_strm1_tmp     ;
  reg [31:0] pe30_lane21_strm0 [0:4095];
  reg [31:0] pe30_lane21_strm0_tmp     ;
  reg [31:0] pe30_lane21_strm1 [0:4095];
  reg [31:0] pe30_lane21_strm1_tmp     ;
  reg [31:0] pe30_lane22_strm0 [0:4095];
  reg [31:0] pe30_lane22_strm0_tmp     ;
  reg [31:0] pe30_lane22_strm1 [0:4095];
  reg [31:0] pe30_lane22_strm1_tmp     ;
  reg [31:0] pe30_lane23_strm0 [0:4095];
  reg [31:0] pe30_lane23_strm0_tmp     ;
  reg [31:0] pe30_lane23_strm1 [0:4095];
  reg [31:0] pe30_lane23_strm1_tmp     ;
  reg [31:0] pe30_lane24_strm0 [0:4095];
  reg [31:0] pe30_lane24_strm0_tmp     ;
  reg [31:0] pe30_lane24_strm1 [0:4095];
  reg [31:0] pe30_lane24_strm1_tmp     ;
  reg [31:0] pe30_lane25_strm0 [0:4095];
  reg [31:0] pe30_lane25_strm0_tmp     ;
  reg [31:0] pe30_lane25_strm1 [0:4095];
  reg [31:0] pe30_lane25_strm1_tmp     ;
  reg [31:0] pe30_lane26_strm0 [0:4095];
  reg [31:0] pe30_lane26_strm0_tmp     ;
  reg [31:0] pe30_lane26_strm1 [0:4095];
  reg [31:0] pe30_lane26_strm1_tmp     ;
  reg [31:0] pe30_lane27_strm0 [0:4095];
  reg [31:0] pe30_lane27_strm0_tmp     ;
  reg [31:0] pe30_lane27_strm1 [0:4095];
  reg [31:0] pe30_lane27_strm1_tmp     ;
  reg [31:0] pe30_lane28_strm0 [0:4095];
  reg [31:0] pe30_lane28_strm0_tmp     ;
  reg [31:0] pe30_lane28_strm1 [0:4095];
  reg [31:0] pe30_lane28_strm1_tmp     ;
  reg [31:0] pe30_lane29_strm0 [0:4095];
  reg [31:0] pe30_lane29_strm0_tmp     ;
  reg [31:0] pe30_lane29_strm1 [0:4095];
  reg [31:0] pe30_lane29_strm1_tmp     ;
  reg [31:0] pe30_lane30_strm0 [0:4095];
  reg [31:0] pe30_lane30_strm0_tmp     ;
  reg [31:0] pe30_lane30_strm1 [0:4095];
  reg [31:0] pe30_lane30_strm1_tmp     ;
  reg [31:0] pe30_lane31_strm0 [0:4095];
  reg [31:0] pe30_lane31_strm0_tmp     ;
  reg [31:0] pe30_lane31_strm1 [0:4095];
  reg [31:0] pe30_lane31_strm1_tmp     ;
  reg [31:0] pe31_lane0_strm0 [0:4095];
  reg [31:0] pe31_lane0_strm0_tmp     ;
  reg [31:0] pe31_lane0_strm1 [0:4095];
  reg [31:0] pe31_lane0_strm1_tmp     ;
  reg [31:0] pe31_lane1_strm0 [0:4095];
  reg [31:0] pe31_lane1_strm0_tmp     ;
  reg [31:0] pe31_lane1_strm1 [0:4095];
  reg [31:0] pe31_lane1_strm1_tmp     ;
  reg [31:0] pe31_lane2_strm0 [0:4095];
  reg [31:0] pe31_lane2_strm0_tmp     ;
  reg [31:0] pe31_lane2_strm1 [0:4095];
  reg [31:0] pe31_lane2_strm1_tmp     ;
  reg [31:0] pe31_lane3_strm0 [0:4095];
  reg [31:0] pe31_lane3_strm0_tmp     ;
  reg [31:0] pe31_lane3_strm1 [0:4095];
  reg [31:0] pe31_lane3_strm1_tmp     ;
  reg [31:0] pe31_lane4_strm0 [0:4095];
  reg [31:0] pe31_lane4_strm0_tmp     ;
  reg [31:0] pe31_lane4_strm1 [0:4095];
  reg [31:0] pe31_lane4_strm1_tmp     ;
  reg [31:0] pe31_lane5_strm0 [0:4095];
  reg [31:0] pe31_lane5_strm0_tmp     ;
  reg [31:0] pe31_lane5_strm1 [0:4095];
  reg [31:0] pe31_lane5_strm1_tmp     ;
  reg [31:0] pe31_lane6_strm0 [0:4095];
  reg [31:0] pe31_lane6_strm0_tmp     ;
  reg [31:0] pe31_lane6_strm1 [0:4095];
  reg [31:0] pe31_lane6_strm1_tmp     ;
  reg [31:0] pe31_lane7_strm0 [0:4095];
  reg [31:0] pe31_lane7_strm0_tmp     ;
  reg [31:0] pe31_lane7_strm1 [0:4095];
  reg [31:0] pe31_lane7_strm1_tmp     ;
  reg [31:0] pe31_lane8_strm0 [0:4095];
  reg [31:0] pe31_lane8_strm0_tmp     ;
  reg [31:0] pe31_lane8_strm1 [0:4095];
  reg [31:0] pe31_lane8_strm1_tmp     ;
  reg [31:0] pe31_lane9_strm0 [0:4095];
  reg [31:0] pe31_lane9_strm0_tmp     ;
  reg [31:0] pe31_lane9_strm1 [0:4095];
  reg [31:0] pe31_lane9_strm1_tmp     ;
  reg [31:0] pe31_lane10_strm0 [0:4095];
  reg [31:0] pe31_lane10_strm0_tmp     ;
  reg [31:0] pe31_lane10_strm1 [0:4095];
  reg [31:0] pe31_lane10_strm1_tmp     ;
  reg [31:0] pe31_lane11_strm0 [0:4095];
  reg [31:0] pe31_lane11_strm0_tmp     ;
  reg [31:0] pe31_lane11_strm1 [0:4095];
  reg [31:0] pe31_lane11_strm1_tmp     ;
  reg [31:0] pe31_lane12_strm0 [0:4095];
  reg [31:0] pe31_lane12_strm0_tmp     ;
  reg [31:0] pe31_lane12_strm1 [0:4095];
  reg [31:0] pe31_lane12_strm1_tmp     ;
  reg [31:0] pe31_lane13_strm0 [0:4095];
  reg [31:0] pe31_lane13_strm0_tmp     ;
  reg [31:0] pe31_lane13_strm1 [0:4095];
  reg [31:0] pe31_lane13_strm1_tmp     ;
  reg [31:0] pe31_lane14_strm0 [0:4095];
  reg [31:0] pe31_lane14_strm0_tmp     ;
  reg [31:0] pe31_lane14_strm1 [0:4095];
  reg [31:0] pe31_lane14_strm1_tmp     ;
  reg [31:0] pe31_lane15_strm0 [0:4095];
  reg [31:0] pe31_lane15_strm0_tmp     ;
  reg [31:0] pe31_lane15_strm1 [0:4095];
  reg [31:0] pe31_lane15_strm1_tmp     ;
  reg [31:0] pe31_lane16_strm0 [0:4095];
  reg [31:0] pe31_lane16_strm0_tmp     ;
  reg [31:0] pe31_lane16_strm1 [0:4095];
  reg [31:0] pe31_lane16_strm1_tmp     ;
  reg [31:0] pe31_lane17_strm0 [0:4095];
  reg [31:0] pe31_lane17_strm0_tmp     ;
  reg [31:0] pe31_lane17_strm1 [0:4095];
  reg [31:0] pe31_lane17_strm1_tmp     ;
  reg [31:0] pe31_lane18_strm0 [0:4095];
  reg [31:0] pe31_lane18_strm0_tmp     ;
  reg [31:0] pe31_lane18_strm1 [0:4095];
  reg [31:0] pe31_lane18_strm1_tmp     ;
  reg [31:0] pe31_lane19_strm0 [0:4095];
  reg [31:0] pe31_lane19_strm0_tmp     ;
  reg [31:0] pe31_lane19_strm1 [0:4095];
  reg [31:0] pe31_lane19_strm1_tmp     ;
  reg [31:0] pe31_lane20_strm0 [0:4095];
  reg [31:0] pe31_lane20_strm0_tmp     ;
  reg [31:0] pe31_lane20_strm1 [0:4095];
  reg [31:0] pe31_lane20_strm1_tmp     ;
  reg [31:0] pe31_lane21_strm0 [0:4095];
  reg [31:0] pe31_lane21_strm0_tmp     ;
  reg [31:0] pe31_lane21_strm1 [0:4095];
  reg [31:0] pe31_lane21_strm1_tmp     ;
  reg [31:0] pe31_lane22_strm0 [0:4095];
  reg [31:0] pe31_lane22_strm0_tmp     ;
  reg [31:0] pe31_lane22_strm1 [0:4095];
  reg [31:0] pe31_lane22_strm1_tmp     ;
  reg [31:0] pe31_lane23_strm0 [0:4095];
  reg [31:0] pe31_lane23_strm0_tmp     ;
  reg [31:0] pe31_lane23_strm1 [0:4095];
  reg [31:0] pe31_lane23_strm1_tmp     ;
  reg [31:0] pe31_lane24_strm0 [0:4095];
  reg [31:0] pe31_lane24_strm0_tmp     ;
  reg [31:0] pe31_lane24_strm1 [0:4095];
  reg [31:0] pe31_lane24_strm1_tmp     ;
  reg [31:0] pe31_lane25_strm0 [0:4095];
  reg [31:0] pe31_lane25_strm0_tmp     ;
  reg [31:0] pe31_lane25_strm1 [0:4095];
  reg [31:0] pe31_lane25_strm1_tmp     ;
  reg [31:0] pe31_lane26_strm0 [0:4095];
  reg [31:0] pe31_lane26_strm0_tmp     ;
  reg [31:0] pe31_lane26_strm1 [0:4095];
  reg [31:0] pe31_lane26_strm1_tmp     ;
  reg [31:0] pe31_lane27_strm0 [0:4095];
  reg [31:0] pe31_lane27_strm0_tmp     ;
  reg [31:0] pe31_lane27_strm1 [0:4095];
  reg [31:0] pe31_lane27_strm1_tmp     ;
  reg [31:0] pe31_lane28_strm0 [0:4095];
  reg [31:0] pe31_lane28_strm0_tmp     ;
  reg [31:0] pe31_lane28_strm1 [0:4095];
  reg [31:0] pe31_lane28_strm1_tmp     ;
  reg [31:0] pe31_lane29_strm0 [0:4095];
  reg [31:0] pe31_lane29_strm0_tmp     ;
  reg [31:0] pe31_lane29_strm1 [0:4095];
  reg [31:0] pe31_lane29_strm1_tmp     ;
  reg [31:0] pe31_lane30_strm0 [0:4095];
  reg [31:0] pe31_lane30_strm0_tmp     ;
  reg [31:0] pe31_lane30_strm1 [0:4095];
  reg [31:0] pe31_lane30_strm1_tmp     ;
  reg [31:0] pe31_lane31_strm0 [0:4095];
  reg [31:0] pe31_lane31_strm0_tmp     ;
  reg [31:0] pe31_lane31_strm1 [0:4095];
  reg [31:0] pe31_lane31_strm1_tmp     ;
  reg [31:0] pe32_lane0_strm0 [0:4095];
  reg [31:0] pe32_lane0_strm0_tmp     ;
  reg [31:0] pe32_lane0_strm1 [0:4095];
  reg [31:0] pe32_lane0_strm1_tmp     ;
  reg [31:0] pe32_lane1_strm0 [0:4095];
  reg [31:0] pe32_lane1_strm0_tmp     ;
  reg [31:0] pe32_lane1_strm1 [0:4095];
  reg [31:0] pe32_lane1_strm1_tmp     ;
  reg [31:0] pe32_lane2_strm0 [0:4095];
  reg [31:0] pe32_lane2_strm0_tmp     ;
  reg [31:0] pe32_lane2_strm1 [0:4095];
  reg [31:0] pe32_lane2_strm1_tmp     ;
  reg [31:0] pe32_lane3_strm0 [0:4095];
  reg [31:0] pe32_lane3_strm0_tmp     ;
  reg [31:0] pe32_lane3_strm1 [0:4095];
  reg [31:0] pe32_lane3_strm1_tmp     ;
  reg [31:0] pe32_lane4_strm0 [0:4095];
  reg [31:0] pe32_lane4_strm0_tmp     ;
  reg [31:0] pe32_lane4_strm1 [0:4095];
  reg [31:0] pe32_lane4_strm1_tmp     ;
  reg [31:0] pe32_lane5_strm0 [0:4095];
  reg [31:0] pe32_lane5_strm0_tmp     ;
  reg [31:0] pe32_lane5_strm1 [0:4095];
  reg [31:0] pe32_lane5_strm1_tmp     ;
  reg [31:0] pe32_lane6_strm0 [0:4095];
  reg [31:0] pe32_lane6_strm0_tmp     ;
  reg [31:0] pe32_lane6_strm1 [0:4095];
  reg [31:0] pe32_lane6_strm1_tmp     ;
  reg [31:0] pe32_lane7_strm0 [0:4095];
  reg [31:0] pe32_lane7_strm0_tmp     ;
  reg [31:0] pe32_lane7_strm1 [0:4095];
  reg [31:0] pe32_lane7_strm1_tmp     ;
  reg [31:0] pe32_lane8_strm0 [0:4095];
  reg [31:0] pe32_lane8_strm0_tmp     ;
  reg [31:0] pe32_lane8_strm1 [0:4095];
  reg [31:0] pe32_lane8_strm1_tmp     ;
  reg [31:0] pe32_lane9_strm0 [0:4095];
  reg [31:0] pe32_lane9_strm0_tmp     ;
  reg [31:0] pe32_lane9_strm1 [0:4095];
  reg [31:0] pe32_lane9_strm1_tmp     ;
  reg [31:0] pe32_lane10_strm0 [0:4095];
  reg [31:0] pe32_lane10_strm0_tmp     ;
  reg [31:0] pe32_lane10_strm1 [0:4095];
  reg [31:0] pe32_lane10_strm1_tmp     ;
  reg [31:0] pe32_lane11_strm0 [0:4095];
  reg [31:0] pe32_lane11_strm0_tmp     ;
  reg [31:0] pe32_lane11_strm1 [0:4095];
  reg [31:0] pe32_lane11_strm1_tmp     ;
  reg [31:0] pe32_lane12_strm0 [0:4095];
  reg [31:0] pe32_lane12_strm0_tmp     ;
  reg [31:0] pe32_lane12_strm1 [0:4095];
  reg [31:0] pe32_lane12_strm1_tmp     ;
  reg [31:0] pe32_lane13_strm0 [0:4095];
  reg [31:0] pe32_lane13_strm0_tmp     ;
  reg [31:0] pe32_lane13_strm1 [0:4095];
  reg [31:0] pe32_lane13_strm1_tmp     ;
  reg [31:0] pe32_lane14_strm0 [0:4095];
  reg [31:0] pe32_lane14_strm0_tmp     ;
  reg [31:0] pe32_lane14_strm1 [0:4095];
  reg [31:0] pe32_lane14_strm1_tmp     ;
  reg [31:0] pe32_lane15_strm0 [0:4095];
  reg [31:0] pe32_lane15_strm0_tmp     ;
  reg [31:0] pe32_lane15_strm1 [0:4095];
  reg [31:0] pe32_lane15_strm1_tmp     ;
  reg [31:0] pe32_lane16_strm0 [0:4095];
  reg [31:0] pe32_lane16_strm0_tmp     ;
  reg [31:0] pe32_lane16_strm1 [0:4095];
  reg [31:0] pe32_lane16_strm1_tmp     ;
  reg [31:0] pe32_lane17_strm0 [0:4095];
  reg [31:0] pe32_lane17_strm0_tmp     ;
  reg [31:0] pe32_lane17_strm1 [0:4095];
  reg [31:0] pe32_lane17_strm1_tmp     ;
  reg [31:0] pe32_lane18_strm0 [0:4095];
  reg [31:0] pe32_lane18_strm0_tmp     ;
  reg [31:0] pe32_lane18_strm1 [0:4095];
  reg [31:0] pe32_lane18_strm1_tmp     ;
  reg [31:0] pe32_lane19_strm0 [0:4095];
  reg [31:0] pe32_lane19_strm0_tmp     ;
  reg [31:0] pe32_lane19_strm1 [0:4095];
  reg [31:0] pe32_lane19_strm1_tmp     ;
  reg [31:0] pe32_lane20_strm0 [0:4095];
  reg [31:0] pe32_lane20_strm0_tmp     ;
  reg [31:0] pe32_lane20_strm1 [0:4095];
  reg [31:0] pe32_lane20_strm1_tmp     ;
  reg [31:0] pe32_lane21_strm0 [0:4095];
  reg [31:0] pe32_lane21_strm0_tmp     ;
  reg [31:0] pe32_lane21_strm1 [0:4095];
  reg [31:0] pe32_lane21_strm1_tmp     ;
  reg [31:0] pe32_lane22_strm0 [0:4095];
  reg [31:0] pe32_lane22_strm0_tmp     ;
  reg [31:0] pe32_lane22_strm1 [0:4095];
  reg [31:0] pe32_lane22_strm1_tmp     ;
  reg [31:0] pe32_lane23_strm0 [0:4095];
  reg [31:0] pe32_lane23_strm0_tmp     ;
  reg [31:0] pe32_lane23_strm1 [0:4095];
  reg [31:0] pe32_lane23_strm1_tmp     ;
  reg [31:0] pe32_lane24_strm0 [0:4095];
  reg [31:0] pe32_lane24_strm0_tmp     ;
  reg [31:0] pe32_lane24_strm1 [0:4095];
  reg [31:0] pe32_lane24_strm1_tmp     ;
  reg [31:0] pe32_lane25_strm0 [0:4095];
  reg [31:0] pe32_lane25_strm0_tmp     ;
  reg [31:0] pe32_lane25_strm1 [0:4095];
  reg [31:0] pe32_lane25_strm1_tmp     ;
  reg [31:0] pe32_lane26_strm0 [0:4095];
  reg [31:0] pe32_lane26_strm0_tmp     ;
  reg [31:0] pe32_lane26_strm1 [0:4095];
  reg [31:0] pe32_lane26_strm1_tmp     ;
  reg [31:0] pe32_lane27_strm0 [0:4095];
  reg [31:0] pe32_lane27_strm0_tmp     ;
  reg [31:0] pe32_lane27_strm1 [0:4095];
  reg [31:0] pe32_lane27_strm1_tmp     ;
  reg [31:0] pe32_lane28_strm0 [0:4095];
  reg [31:0] pe32_lane28_strm0_tmp     ;
  reg [31:0] pe32_lane28_strm1 [0:4095];
  reg [31:0] pe32_lane28_strm1_tmp     ;
  reg [31:0] pe32_lane29_strm0 [0:4095];
  reg [31:0] pe32_lane29_strm0_tmp     ;
  reg [31:0] pe32_lane29_strm1 [0:4095];
  reg [31:0] pe32_lane29_strm1_tmp     ;
  reg [31:0] pe32_lane30_strm0 [0:4095];
  reg [31:0] pe32_lane30_strm0_tmp     ;
  reg [31:0] pe32_lane30_strm1 [0:4095];
  reg [31:0] pe32_lane30_strm1_tmp     ;
  reg [31:0] pe32_lane31_strm0 [0:4095];
  reg [31:0] pe32_lane31_strm0_tmp     ;
  reg [31:0] pe32_lane31_strm1 [0:4095];
  reg [31:0] pe32_lane31_strm1_tmp     ;
  reg [31:0] pe33_lane0_strm0 [0:4095];
  reg [31:0] pe33_lane0_strm0_tmp     ;
  reg [31:0] pe33_lane0_strm1 [0:4095];
  reg [31:0] pe33_lane0_strm1_tmp     ;
  reg [31:0] pe33_lane1_strm0 [0:4095];
  reg [31:0] pe33_lane1_strm0_tmp     ;
  reg [31:0] pe33_lane1_strm1 [0:4095];
  reg [31:0] pe33_lane1_strm1_tmp     ;
  reg [31:0] pe33_lane2_strm0 [0:4095];
  reg [31:0] pe33_lane2_strm0_tmp     ;
  reg [31:0] pe33_lane2_strm1 [0:4095];
  reg [31:0] pe33_lane2_strm1_tmp     ;
  reg [31:0] pe33_lane3_strm0 [0:4095];
  reg [31:0] pe33_lane3_strm0_tmp     ;
  reg [31:0] pe33_lane3_strm1 [0:4095];
  reg [31:0] pe33_lane3_strm1_tmp     ;
  reg [31:0] pe33_lane4_strm0 [0:4095];
  reg [31:0] pe33_lane4_strm0_tmp     ;
  reg [31:0] pe33_lane4_strm1 [0:4095];
  reg [31:0] pe33_lane4_strm1_tmp     ;
  reg [31:0] pe33_lane5_strm0 [0:4095];
  reg [31:0] pe33_lane5_strm0_tmp     ;
  reg [31:0] pe33_lane5_strm1 [0:4095];
  reg [31:0] pe33_lane5_strm1_tmp     ;
  reg [31:0] pe33_lane6_strm0 [0:4095];
  reg [31:0] pe33_lane6_strm0_tmp     ;
  reg [31:0] pe33_lane6_strm1 [0:4095];
  reg [31:0] pe33_lane6_strm1_tmp     ;
  reg [31:0] pe33_lane7_strm0 [0:4095];
  reg [31:0] pe33_lane7_strm0_tmp     ;
  reg [31:0] pe33_lane7_strm1 [0:4095];
  reg [31:0] pe33_lane7_strm1_tmp     ;
  reg [31:0] pe33_lane8_strm0 [0:4095];
  reg [31:0] pe33_lane8_strm0_tmp     ;
  reg [31:0] pe33_lane8_strm1 [0:4095];
  reg [31:0] pe33_lane8_strm1_tmp     ;
  reg [31:0] pe33_lane9_strm0 [0:4095];
  reg [31:0] pe33_lane9_strm0_tmp     ;
  reg [31:0] pe33_lane9_strm1 [0:4095];
  reg [31:0] pe33_lane9_strm1_tmp     ;
  reg [31:0] pe33_lane10_strm0 [0:4095];
  reg [31:0] pe33_lane10_strm0_tmp     ;
  reg [31:0] pe33_lane10_strm1 [0:4095];
  reg [31:0] pe33_lane10_strm1_tmp     ;
  reg [31:0] pe33_lane11_strm0 [0:4095];
  reg [31:0] pe33_lane11_strm0_tmp     ;
  reg [31:0] pe33_lane11_strm1 [0:4095];
  reg [31:0] pe33_lane11_strm1_tmp     ;
  reg [31:0] pe33_lane12_strm0 [0:4095];
  reg [31:0] pe33_lane12_strm0_tmp     ;
  reg [31:0] pe33_lane12_strm1 [0:4095];
  reg [31:0] pe33_lane12_strm1_tmp     ;
  reg [31:0] pe33_lane13_strm0 [0:4095];
  reg [31:0] pe33_lane13_strm0_tmp     ;
  reg [31:0] pe33_lane13_strm1 [0:4095];
  reg [31:0] pe33_lane13_strm1_tmp     ;
  reg [31:0] pe33_lane14_strm0 [0:4095];
  reg [31:0] pe33_lane14_strm0_tmp     ;
  reg [31:0] pe33_lane14_strm1 [0:4095];
  reg [31:0] pe33_lane14_strm1_tmp     ;
  reg [31:0] pe33_lane15_strm0 [0:4095];
  reg [31:0] pe33_lane15_strm0_tmp     ;
  reg [31:0] pe33_lane15_strm1 [0:4095];
  reg [31:0] pe33_lane15_strm1_tmp     ;
  reg [31:0] pe33_lane16_strm0 [0:4095];
  reg [31:0] pe33_lane16_strm0_tmp     ;
  reg [31:0] pe33_lane16_strm1 [0:4095];
  reg [31:0] pe33_lane16_strm1_tmp     ;
  reg [31:0] pe33_lane17_strm0 [0:4095];
  reg [31:0] pe33_lane17_strm0_tmp     ;
  reg [31:0] pe33_lane17_strm1 [0:4095];
  reg [31:0] pe33_lane17_strm1_tmp     ;
  reg [31:0] pe33_lane18_strm0 [0:4095];
  reg [31:0] pe33_lane18_strm0_tmp     ;
  reg [31:0] pe33_lane18_strm1 [0:4095];
  reg [31:0] pe33_lane18_strm1_tmp     ;
  reg [31:0] pe33_lane19_strm0 [0:4095];
  reg [31:0] pe33_lane19_strm0_tmp     ;
  reg [31:0] pe33_lane19_strm1 [0:4095];
  reg [31:0] pe33_lane19_strm1_tmp     ;
  reg [31:0] pe33_lane20_strm0 [0:4095];
  reg [31:0] pe33_lane20_strm0_tmp     ;
  reg [31:0] pe33_lane20_strm1 [0:4095];
  reg [31:0] pe33_lane20_strm1_tmp     ;
  reg [31:0] pe33_lane21_strm0 [0:4095];
  reg [31:0] pe33_lane21_strm0_tmp     ;
  reg [31:0] pe33_lane21_strm1 [0:4095];
  reg [31:0] pe33_lane21_strm1_tmp     ;
  reg [31:0] pe33_lane22_strm0 [0:4095];
  reg [31:0] pe33_lane22_strm0_tmp     ;
  reg [31:0] pe33_lane22_strm1 [0:4095];
  reg [31:0] pe33_lane22_strm1_tmp     ;
  reg [31:0] pe33_lane23_strm0 [0:4095];
  reg [31:0] pe33_lane23_strm0_tmp     ;
  reg [31:0] pe33_lane23_strm1 [0:4095];
  reg [31:0] pe33_lane23_strm1_tmp     ;
  reg [31:0] pe33_lane24_strm0 [0:4095];
  reg [31:0] pe33_lane24_strm0_tmp     ;
  reg [31:0] pe33_lane24_strm1 [0:4095];
  reg [31:0] pe33_lane24_strm1_tmp     ;
  reg [31:0] pe33_lane25_strm0 [0:4095];
  reg [31:0] pe33_lane25_strm0_tmp     ;
  reg [31:0] pe33_lane25_strm1 [0:4095];
  reg [31:0] pe33_lane25_strm1_tmp     ;
  reg [31:0] pe33_lane26_strm0 [0:4095];
  reg [31:0] pe33_lane26_strm0_tmp     ;
  reg [31:0] pe33_lane26_strm1 [0:4095];
  reg [31:0] pe33_lane26_strm1_tmp     ;
  reg [31:0] pe33_lane27_strm0 [0:4095];
  reg [31:0] pe33_lane27_strm0_tmp     ;
  reg [31:0] pe33_lane27_strm1 [0:4095];
  reg [31:0] pe33_lane27_strm1_tmp     ;
  reg [31:0] pe33_lane28_strm0 [0:4095];
  reg [31:0] pe33_lane28_strm0_tmp     ;
  reg [31:0] pe33_lane28_strm1 [0:4095];
  reg [31:0] pe33_lane28_strm1_tmp     ;
  reg [31:0] pe33_lane29_strm0 [0:4095];
  reg [31:0] pe33_lane29_strm0_tmp     ;
  reg [31:0] pe33_lane29_strm1 [0:4095];
  reg [31:0] pe33_lane29_strm1_tmp     ;
  reg [31:0] pe33_lane30_strm0 [0:4095];
  reg [31:0] pe33_lane30_strm0_tmp     ;
  reg [31:0] pe33_lane30_strm1 [0:4095];
  reg [31:0] pe33_lane30_strm1_tmp     ;
  reg [31:0] pe33_lane31_strm0 [0:4095];
  reg [31:0] pe33_lane31_strm0_tmp     ;
  reg [31:0] pe33_lane31_strm1 [0:4095];
  reg [31:0] pe33_lane31_strm1_tmp     ;
  reg [31:0] pe34_lane0_strm0 [0:4095];
  reg [31:0] pe34_lane0_strm0_tmp     ;
  reg [31:0] pe34_lane0_strm1 [0:4095];
  reg [31:0] pe34_lane0_strm1_tmp     ;
  reg [31:0] pe34_lane1_strm0 [0:4095];
  reg [31:0] pe34_lane1_strm0_tmp     ;
  reg [31:0] pe34_lane1_strm1 [0:4095];
  reg [31:0] pe34_lane1_strm1_tmp     ;
  reg [31:0] pe34_lane2_strm0 [0:4095];
  reg [31:0] pe34_lane2_strm0_tmp     ;
  reg [31:0] pe34_lane2_strm1 [0:4095];
  reg [31:0] pe34_lane2_strm1_tmp     ;
  reg [31:0] pe34_lane3_strm0 [0:4095];
  reg [31:0] pe34_lane3_strm0_tmp     ;
  reg [31:0] pe34_lane3_strm1 [0:4095];
  reg [31:0] pe34_lane3_strm1_tmp     ;
  reg [31:0] pe34_lane4_strm0 [0:4095];
  reg [31:0] pe34_lane4_strm0_tmp     ;
  reg [31:0] pe34_lane4_strm1 [0:4095];
  reg [31:0] pe34_lane4_strm1_tmp     ;
  reg [31:0] pe34_lane5_strm0 [0:4095];
  reg [31:0] pe34_lane5_strm0_tmp     ;
  reg [31:0] pe34_lane5_strm1 [0:4095];
  reg [31:0] pe34_lane5_strm1_tmp     ;
  reg [31:0] pe34_lane6_strm0 [0:4095];
  reg [31:0] pe34_lane6_strm0_tmp     ;
  reg [31:0] pe34_lane6_strm1 [0:4095];
  reg [31:0] pe34_lane6_strm1_tmp     ;
  reg [31:0] pe34_lane7_strm0 [0:4095];
  reg [31:0] pe34_lane7_strm0_tmp     ;
  reg [31:0] pe34_lane7_strm1 [0:4095];
  reg [31:0] pe34_lane7_strm1_tmp     ;
  reg [31:0] pe34_lane8_strm0 [0:4095];
  reg [31:0] pe34_lane8_strm0_tmp     ;
  reg [31:0] pe34_lane8_strm1 [0:4095];
  reg [31:0] pe34_lane8_strm1_tmp     ;
  reg [31:0] pe34_lane9_strm0 [0:4095];
  reg [31:0] pe34_lane9_strm0_tmp     ;
  reg [31:0] pe34_lane9_strm1 [0:4095];
  reg [31:0] pe34_lane9_strm1_tmp     ;
  reg [31:0] pe34_lane10_strm0 [0:4095];
  reg [31:0] pe34_lane10_strm0_tmp     ;
  reg [31:0] pe34_lane10_strm1 [0:4095];
  reg [31:0] pe34_lane10_strm1_tmp     ;
  reg [31:0] pe34_lane11_strm0 [0:4095];
  reg [31:0] pe34_lane11_strm0_tmp     ;
  reg [31:0] pe34_lane11_strm1 [0:4095];
  reg [31:0] pe34_lane11_strm1_tmp     ;
  reg [31:0] pe34_lane12_strm0 [0:4095];
  reg [31:0] pe34_lane12_strm0_tmp     ;
  reg [31:0] pe34_lane12_strm1 [0:4095];
  reg [31:0] pe34_lane12_strm1_tmp     ;
  reg [31:0] pe34_lane13_strm0 [0:4095];
  reg [31:0] pe34_lane13_strm0_tmp     ;
  reg [31:0] pe34_lane13_strm1 [0:4095];
  reg [31:0] pe34_lane13_strm1_tmp     ;
  reg [31:0] pe34_lane14_strm0 [0:4095];
  reg [31:0] pe34_lane14_strm0_tmp     ;
  reg [31:0] pe34_lane14_strm1 [0:4095];
  reg [31:0] pe34_lane14_strm1_tmp     ;
  reg [31:0] pe34_lane15_strm0 [0:4095];
  reg [31:0] pe34_lane15_strm0_tmp     ;
  reg [31:0] pe34_lane15_strm1 [0:4095];
  reg [31:0] pe34_lane15_strm1_tmp     ;
  reg [31:0] pe34_lane16_strm0 [0:4095];
  reg [31:0] pe34_lane16_strm0_tmp     ;
  reg [31:0] pe34_lane16_strm1 [0:4095];
  reg [31:0] pe34_lane16_strm1_tmp     ;
  reg [31:0] pe34_lane17_strm0 [0:4095];
  reg [31:0] pe34_lane17_strm0_tmp     ;
  reg [31:0] pe34_lane17_strm1 [0:4095];
  reg [31:0] pe34_lane17_strm1_tmp     ;
  reg [31:0] pe34_lane18_strm0 [0:4095];
  reg [31:0] pe34_lane18_strm0_tmp     ;
  reg [31:0] pe34_lane18_strm1 [0:4095];
  reg [31:0] pe34_lane18_strm1_tmp     ;
  reg [31:0] pe34_lane19_strm0 [0:4095];
  reg [31:0] pe34_lane19_strm0_tmp     ;
  reg [31:0] pe34_lane19_strm1 [0:4095];
  reg [31:0] pe34_lane19_strm1_tmp     ;
  reg [31:0] pe34_lane20_strm0 [0:4095];
  reg [31:0] pe34_lane20_strm0_tmp     ;
  reg [31:0] pe34_lane20_strm1 [0:4095];
  reg [31:0] pe34_lane20_strm1_tmp     ;
  reg [31:0] pe34_lane21_strm0 [0:4095];
  reg [31:0] pe34_lane21_strm0_tmp     ;
  reg [31:0] pe34_lane21_strm1 [0:4095];
  reg [31:0] pe34_lane21_strm1_tmp     ;
  reg [31:0] pe34_lane22_strm0 [0:4095];
  reg [31:0] pe34_lane22_strm0_tmp     ;
  reg [31:0] pe34_lane22_strm1 [0:4095];
  reg [31:0] pe34_lane22_strm1_tmp     ;
  reg [31:0] pe34_lane23_strm0 [0:4095];
  reg [31:0] pe34_lane23_strm0_tmp     ;
  reg [31:0] pe34_lane23_strm1 [0:4095];
  reg [31:0] pe34_lane23_strm1_tmp     ;
  reg [31:0] pe34_lane24_strm0 [0:4095];
  reg [31:0] pe34_lane24_strm0_tmp     ;
  reg [31:0] pe34_lane24_strm1 [0:4095];
  reg [31:0] pe34_lane24_strm1_tmp     ;
  reg [31:0] pe34_lane25_strm0 [0:4095];
  reg [31:0] pe34_lane25_strm0_tmp     ;
  reg [31:0] pe34_lane25_strm1 [0:4095];
  reg [31:0] pe34_lane25_strm1_tmp     ;
  reg [31:0] pe34_lane26_strm0 [0:4095];
  reg [31:0] pe34_lane26_strm0_tmp     ;
  reg [31:0] pe34_lane26_strm1 [0:4095];
  reg [31:0] pe34_lane26_strm1_tmp     ;
  reg [31:0] pe34_lane27_strm0 [0:4095];
  reg [31:0] pe34_lane27_strm0_tmp     ;
  reg [31:0] pe34_lane27_strm1 [0:4095];
  reg [31:0] pe34_lane27_strm1_tmp     ;
  reg [31:0] pe34_lane28_strm0 [0:4095];
  reg [31:0] pe34_lane28_strm0_tmp     ;
  reg [31:0] pe34_lane28_strm1 [0:4095];
  reg [31:0] pe34_lane28_strm1_tmp     ;
  reg [31:0] pe34_lane29_strm0 [0:4095];
  reg [31:0] pe34_lane29_strm0_tmp     ;
  reg [31:0] pe34_lane29_strm1 [0:4095];
  reg [31:0] pe34_lane29_strm1_tmp     ;
  reg [31:0] pe34_lane30_strm0 [0:4095];
  reg [31:0] pe34_lane30_strm0_tmp     ;
  reg [31:0] pe34_lane30_strm1 [0:4095];
  reg [31:0] pe34_lane30_strm1_tmp     ;
  reg [31:0] pe34_lane31_strm0 [0:4095];
  reg [31:0] pe34_lane31_strm0_tmp     ;
  reg [31:0] pe34_lane31_strm1 [0:4095];
  reg [31:0] pe34_lane31_strm1_tmp     ;
  reg [31:0] pe35_lane0_strm0 [0:4095];
  reg [31:0] pe35_lane0_strm0_tmp     ;
  reg [31:0] pe35_lane0_strm1 [0:4095];
  reg [31:0] pe35_lane0_strm1_tmp     ;
  reg [31:0] pe35_lane1_strm0 [0:4095];
  reg [31:0] pe35_lane1_strm0_tmp     ;
  reg [31:0] pe35_lane1_strm1 [0:4095];
  reg [31:0] pe35_lane1_strm1_tmp     ;
  reg [31:0] pe35_lane2_strm0 [0:4095];
  reg [31:0] pe35_lane2_strm0_tmp     ;
  reg [31:0] pe35_lane2_strm1 [0:4095];
  reg [31:0] pe35_lane2_strm1_tmp     ;
  reg [31:0] pe35_lane3_strm0 [0:4095];
  reg [31:0] pe35_lane3_strm0_tmp     ;
  reg [31:0] pe35_lane3_strm1 [0:4095];
  reg [31:0] pe35_lane3_strm1_tmp     ;
  reg [31:0] pe35_lane4_strm0 [0:4095];
  reg [31:0] pe35_lane4_strm0_tmp     ;
  reg [31:0] pe35_lane4_strm1 [0:4095];
  reg [31:0] pe35_lane4_strm1_tmp     ;
  reg [31:0] pe35_lane5_strm0 [0:4095];
  reg [31:0] pe35_lane5_strm0_tmp     ;
  reg [31:0] pe35_lane5_strm1 [0:4095];
  reg [31:0] pe35_lane5_strm1_tmp     ;
  reg [31:0] pe35_lane6_strm0 [0:4095];
  reg [31:0] pe35_lane6_strm0_tmp     ;
  reg [31:0] pe35_lane6_strm1 [0:4095];
  reg [31:0] pe35_lane6_strm1_tmp     ;
  reg [31:0] pe35_lane7_strm0 [0:4095];
  reg [31:0] pe35_lane7_strm0_tmp     ;
  reg [31:0] pe35_lane7_strm1 [0:4095];
  reg [31:0] pe35_lane7_strm1_tmp     ;
  reg [31:0] pe35_lane8_strm0 [0:4095];
  reg [31:0] pe35_lane8_strm0_tmp     ;
  reg [31:0] pe35_lane8_strm1 [0:4095];
  reg [31:0] pe35_lane8_strm1_tmp     ;
  reg [31:0] pe35_lane9_strm0 [0:4095];
  reg [31:0] pe35_lane9_strm0_tmp     ;
  reg [31:0] pe35_lane9_strm1 [0:4095];
  reg [31:0] pe35_lane9_strm1_tmp     ;
  reg [31:0] pe35_lane10_strm0 [0:4095];
  reg [31:0] pe35_lane10_strm0_tmp     ;
  reg [31:0] pe35_lane10_strm1 [0:4095];
  reg [31:0] pe35_lane10_strm1_tmp     ;
  reg [31:0] pe35_lane11_strm0 [0:4095];
  reg [31:0] pe35_lane11_strm0_tmp     ;
  reg [31:0] pe35_lane11_strm1 [0:4095];
  reg [31:0] pe35_lane11_strm1_tmp     ;
  reg [31:0] pe35_lane12_strm0 [0:4095];
  reg [31:0] pe35_lane12_strm0_tmp     ;
  reg [31:0] pe35_lane12_strm1 [0:4095];
  reg [31:0] pe35_lane12_strm1_tmp     ;
  reg [31:0] pe35_lane13_strm0 [0:4095];
  reg [31:0] pe35_lane13_strm0_tmp     ;
  reg [31:0] pe35_lane13_strm1 [0:4095];
  reg [31:0] pe35_lane13_strm1_tmp     ;
  reg [31:0] pe35_lane14_strm0 [0:4095];
  reg [31:0] pe35_lane14_strm0_tmp     ;
  reg [31:0] pe35_lane14_strm1 [0:4095];
  reg [31:0] pe35_lane14_strm1_tmp     ;
  reg [31:0] pe35_lane15_strm0 [0:4095];
  reg [31:0] pe35_lane15_strm0_tmp     ;
  reg [31:0] pe35_lane15_strm1 [0:4095];
  reg [31:0] pe35_lane15_strm1_tmp     ;
  reg [31:0] pe35_lane16_strm0 [0:4095];
  reg [31:0] pe35_lane16_strm0_tmp     ;
  reg [31:0] pe35_lane16_strm1 [0:4095];
  reg [31:0] pe35_lane16_strm1_tmp     ;
  reg [31:0] pe35_lane17_strm0 [0:4095];
  reg [31:0] pe35_lane17_strm0_tmp     ;
  reg [31:0] pe35_lane17_strm1 [0:4095];
  reg [31:0] pe35_lane17_strm1_tmp     ;
  reg [31:0] pe35_lane18_strm0 [0:4095];
  reg [31:0] pe35_lane18_strm0_tmp     ;
  reg [31:0] pe35_lane18_strm1 [0:4095];
  reg [31:0] pe35_lane18_strm1_tmp     ;
  reg [31:0] pe35_lane19_strm0 [0:4095];
  reg [31:0] pe35_lane19_strm0_tmp     ;
  reg [31:0] pe35_lane19_strm1 [0:4095];
  reg [31:0] pe35_lane19_strm1_tmp     ;
  reg [31:0] pe35_lane20_strm0 [0:4095];
  reg [31:0] pe35_lane20_strm0_tmp     ;
  reg [31:0] pe35_lane20_strm1 [0:4095];
  reg [31:0] pe35_lane20_strm1_tmp     ;
  reg [31:0] pe35_lane21_strm0 [0:4095];
  reg [31:0] pe35_lane21_strm0_tmp     ;
  reg [31:0] pe35_lane21_strm1 [0:4095];
  reg [31:0] pe35_lane21_strm1_tmp     ;
  reg [31:0] pe35_lane22_strm0 [0:4095];
  reg [31:0] pe35_lane22_strm0_tmp     ;
  reg [31:0] pe35_lane22_strm1 [0:4095];
  reg [31:0] pe35_lane22_strm1_tmp     ;
  reg [31:0] pe35_lane23_strm0 [0:4095];
  reg [31:0] pe35_lane23_strm0_tmp     ;
  reg [31:0] pe35_lane23_strm1 [0:4095];
  reg [31:0] pe35_lane23_strm1_tmp     ;
  reg [31:0] pe35_lane24_strm0 [0:4095];
  reg [31:0] pe35_lane24_strm0_tmp     ;
  reg [31:0] pe35_lane24_strm1 [0:4095];
  reg [31:0] pe35_lane24_strm1_tmp     ;
  reg [31:0] pe35_lane25_strm0 [0:4095];
  reg [31:0] pe35_lane25_strm0_tmp     ;
  reg [31:0] pe35_lane25_strm1 [0:4095];
  reg [31:0] pe35_lane25_strm1_tmp     ;
  reg [31:0] pe35_lane26_strm0 [0:4095];
  reg [31:0] pe35_lane26_strm0_tmp     ;
  reg [31:0] pe35_lane26_strm1 [0:4095];
  reg [31:0] pe35_lane26_strm1_tmp     ;
  reg [31:0] pe35_lane27_strm0 [0:4095];
  reg [31:0] pe35_lane27_strm0_tmp     ;
  reg [31:0] pe35_lane27_strm1 [0:4095];
  reg [31:0] pe35_lane27_strm1_tmp     ;
  reg [31:0] pe35_lane28_strm0 [0:4095];
  reg [31:0] pe35_lane28_strm0_tmp     ;
  reg [31:0] pe35_lane28_strm1 [0:4095];
  reg [31:0] pe35_lane28_strm1_tmp     ;
  reg [31:0] pe35_lane29_strm0 [0:4095];
  reg [31:0] pe35_lane29_strm0_tmp     ;
  reg [31:0] pe35_lane29_strm1 [0:4095];
  reg [31:0] pe35_lane29_strm1_tmp     ;
  reg [31:0] pe35_lane30_strm0 [0:4095];
  reg [31:0] pe35_lane30_strm0_tmp     ;
  reg [31:0] pe35_lane30_strm1 [0:4095];
  reg [31:0] pe35_lane30_strm1_tmp     ;
  reg [31:0] pe35_lane31_strm0 [0:4095];
  reg [31:0] pe35_lane31_strm0_tmp     ;
  reg [31:0] pe35_lane31_strm1 [0:4095];
  reg [31:0] pe35_lane31_strm1_tmp     ;
  reg [31:0] pe36_lane0_strm0 [0:4095];
  reg [31:0] pe36_lane0_strm0_tmp     ;
  reg [31:0] pe36_lane0_strm1 [0:4095];
  reg [31:0] pe36_lane0_strm1_tmp     ;
  reg [31:0] pe36_lane1_strm0 [0:4095];
  reg [31:0] pe36_lane1_strm0_tmp     ;
  reg [31:0] pe36_lane1_strm1 [0:4095];
  reg [31:0] pe36_lane1_strm1_tmp     ;
  reg [31:0] pe36_lane2_strm0 [0:4095];
  reg [31:0] pe36_lane2_strm0_tmp     ;
  reg [31:0] pe36_lane2_strm1 [0:4095];
  reg [31:0] pe36_lane2_strm1_tmp     ;
  reg [31:0] pe36_lane3_strm0 [0:4095];
  reg [31:0] pe36_lane3_strm0_tmp     ;
  reg [31:0] pe36_lane3_strm1 [0:4095];
  reg [31:0] pe36_lane3_strm1_tmp     ;
  reg [31:0] pe36_lane4_strm0 [0:4095];
  reg [31:0] pe36_lane4_strm0_tmp     ;
  reg [31:0] pe36_lane4_strm1 [0:4095];
  reg [31:0] pe36_lane4_strm1_tmp     ;
  reg [31:0] pe36_lane5_strm0 [0:4095];
  reg [31:0] pe36_lane5_strm0_tmp     ;
  reg [31:0] pe36_lane5_strm1 [0:4095];
  reg [31:0] pe36_lane5_strm1_tmp     ;
  reg [31:0] pe36_lane6_strm0 [0:4095];
  reg [31:0] pe36_lane6_strm0_tmp     ;
  reg [31:0] pe36_lane6_strm1 [0:4095];
  reg [31:0] pe36_lane6_strm1_tmp     ;
  reg [31:0] pe36_lane7_strm0 [0:4095];
  reg [31:0] pe36_lane7_strm0_tmp     ;
  reg [31:0] pe36_lane7_strm1 [0:4095];
  reg [31:0] pe36_lane7_strm1_tmp     ;
  reg [31:0] pe36_lane8_strm0 [0:4095];
  reg [31:0] pe36_lane8_strm0_tmp     ;
  reg [31:0] pe36_lane8_strm1 [0:4095];
  reg [31:0] pe36_lane8_strm1_tmp     ;
  reg [31:0] pe36_lane9_strm0 [0:4095];
  reg [31:0] pe36_lane9_strm0_tmp     ;
  reg [31:0] pe36_lane9_strm1 [0:4095];
  reg [31:0] pe36_lane9_strm1_tmp     ;
  reg [31:0] pe36_lane10_strm0 [0:4095];
  reg [31:0] pe36_lane10_strm0_tmp     ;
  reg [31:0] pe36_lane10_strm1 [0:4095];
  reg [31:0] pe36_lane10_strm1_tmp     ;
  reg [31:0] pe36_lane11_strm0 [0:4095];
  reg [31:0] pe36_lane11_strm0_tmp     ;
  reg [31:0] pe36_lane11_strm1 [0:4095];
  reg [31:0] pe36_lane11_strm1_tmp     ;
  reg [31:0] pe36_lane12_strm0 [0:4095];
  reg [31:0] pe36_lane12_strm0_tmp     ;
  reg [31:0] pe36_lane12_strm1 [0:4095];
  reg [31:0] pe36_lane12_strm1_tmp     ;
  reg [31:0] pe36_lane13_strm0 [0:4095];
  reg [31:0] pe36_lane13_strm0_tmp     ;
  reg [31:0] pe36_lane13_strm1 [0:4095];
  reg [31:0] pe36_lane13_strm1_tmp     ;
  reg [31:0] pe36_lane14_strm0 [0:4095];
  reg [31:0] pe36_lane14_strm0_tmp     ;
  reg [31:0] pe36_lane14_strm1 [0:4095];
  reg [31:0] pe36_lane14_strm1_tmp     ;
  reg [31:0] pe36_lane15_strm0 [0:4095];
  reg [31:0] pe36_lane15_strm0_tmp     ;
  reg [31:0] pe36_lane15_strm1 [0:4095];
  reg [31:0] pe36_lane15_strm1_tmp     ;
  reg [31:0] pe36_lane16_strm0 [0:4095];
  reg [31:0] pe36_lane16_strm0_tmp     ;
  reg [31:0] pe36_lane16_strm1 [0:4095];
  reg [31:0] pe36_lane16_strm1_tmp     ;
  reg [31:0] pe36_lane17_strm0 [0:4095];
  reg [31:0] pe36_lane17_strm0_tmp     ;
  reg [31:0] pe36_lane17_strm1 [0:4095];
  reg [31:0] pe36_lane17_strm1_tmp     ;
  reg [31:0] pe36_lane18_strm0 [0:4095];
  reg [31:0] pe36_lane18_strm0_tmp     ;
  reg [31:0] pe36_lane18_strm1 [0:4095];
  reg [31:0] pe36_lane18_strm1_tmp     ;
  reg [31:0] pe36_lane19_strm0 [0:4095];
  reg [31:0] pe36_lane19_strm0_tmp     ;
  reg [31:0] pe36_lane19_strm1 [0:4095];
  reg [31:0] pe36_lane19_strm1_tmp     ;
  reg [31:0] pe36_lane20_strm0 [0:4095];
  reg [31:0] pe36_lane20_strm0_tmp     ;
  reg [31:0] pe36_lane20_strm1 [0:4095];
  reg [31:0] pe36_lane20_strm1_tmp     ;
  reg [31:0] pe36_lane21_strm0 [0:4095];
  reg [31:0] pe36_lane21_strm0_tmp     ;
  reg [31:0] pe36_lane21_strm1 [0:4095];
  reg [31:0] pe36_lane21_strm1_tmp     ;
  reg [31:0] pe36_lane22_strm0 [0:4095];
  reg [31:0] pe36_lane22_strm0_tmp     ;
  reg [31:0] pe36_lane22_strm1 [0:4095];
  reg [31:0] pe36_lane22_strm1_tmp     ;
  reg [31:0] pe36_lane23_strm0 [0:4095];
  reg [31:0] pe36_lane23_strm0_tmp     ;
  reg [31:0] pe36_lane23_strm1 [0:4095];
  reg [31:0] pe36_lane23_strm1_tmp     ;
  reg [31:0] pe36_lane24_strm0 [0:4095];
  reg [31:0] pe36_lane24_strm0_tmp     ;
  reg [31:0] pe36_lane24_strm1 [0:4095];
  reg [31:0] pe36_lane24_strm1_tmp     ;
  reg [31:0] pe36_lane25_strm0 [0:4095];
  reg [31:0] pe36_lane25_strm0_tmp     ;
  reg [31:0] pe36_lane25_strm1 [0:4095];
  reg [31:0] pe36_lane25_strm1_tmp     ;
  reg [31:0] pe36_lane26_strm0 [0:4095];
  reg [31:0] pe36_lane26_strm0_tmp     ;
  reg [31:0] pe36_lane26_strm1 [0:4095];
  reg [31:0] pe36_lane26_strm1_tmp     ;
  reg [31:0] pe36_lane27_strm0 [0:4095];
  reg [31:0] pe36_lane27_strm0_tmp     ;
  reg [31:0] pe36_lane27_strm1 [0:4095];
  reg [31:0] pe36_lane27_strm1_tmp     ;
  reg [31:0] pe36_lane28_strm0 [0:4095];
  reg [31:0] pe36_lane28_strm0_tmp     ;
  reg [31:0] pe36_lane28_strm1 [0:4095];
  reg [31:0] pe36_lane28_strm1_tmp     ;
  reg [31:0] pe36_lane29_strm0 [0:4095];
  reg [31:0] pe36_lane29_strm0_tmp     ;
  reg [31:0] pe36_lane29_strm1 [0:4095];
  reg [31:0] pe36_lane29_strm1_tmp     ;
  reg [31:0] pe36_lane30_strm0 [0:4095];
  reg [31:0] pe36_lane30_strm0_tmp     ;
  reg [31:0] pe36_lane30_strm1 [0:4095];
  reg [31:0] pe36_lane30_strm1_tmp     ;
  reg [31:0] pe36_lane31_strm0 [0:4095];
  reg [31:0] pe36_lane31_strm0_tmp     ;
  reg [31:0] pe36_lane31_strm1 [0:4095];
  reg [31:0] pe36_lane31_strm1_tmp     ;
  reg [31:0] pe37_lane0_strm0 [0:4095];
  reg [31:0] pe37_lane0_strm0_tmp     ;
  reg [31:0] pe37_lane0_strm1 [0:4095];
  reg [31:0] pe37_lane0_strm1_tmp     ;
  reg [31:0] pe37_lane1_strm0 [0:4095];
  reg [31:0] pe37_lane1_strm0_tmp     ;
  reg [31:0] pe37_lane1_strm1 [0:4095];
  reg [31:0] pe37_lane1_strm1_tmp     ;
  reg [31:0] pe37_lane2_strm0 [0:4095];
  reg [31:0] pe37_lane2_strm0_tmp     ;
  reg [31:0] pe37_lane2_strm1 [0:4095];
  reg [31:0] pe37_lane2_strm1_tmp     ;
  reg [31:0] pe37_lane3_strm0 [0:4095];
  reg [31:0] pe37_lane3_strm0_tmp     ;
  reg [31:0] pe37_lane3_strm1 [0:4095];
  reg [31:0] pe37_lane3_strm1_tmp     ;
  reg [31:0] pe37_lane4_strm0 [0:4095];
  reg [31:0] pe37_lane4_strm0_tmp     ;
  reg [31:0] pe37_lane4_strm1 [0:4095];
  reg [31:0] pe37_lane4_strm1_tmp     ;
  reg [31:0] pe37_lane5_strm0 [0:4095];
  reg [31:0] pe37_lane5_strm0_tmp     ;
  reg [31:0] pe37_lane5_strm1 [0:4095];
  reg [31:0] pe37_lane5_strm1_tmp     ;
  reg [31:0] pe37_lane6_strm0 [0:4095];
  reg [31:0] pe37_lane6_strm0_tmp     ;
  reg [31:0] pe37_lane6_strm1 [0:4095];
  reg [31:0] pe37_lane6_strm1_tmp     ;
  reg [31:0] pe37_lane7_strm0 [0:4095];
  reg [31:0] pe37_lane7_strm0_tmp     ;
  reg [31:0] pe37_lane7_strm1 [0:4095];
  reg [31:0] pe37_lane7_strm1_tmp     ;
  reg [31:0] pe37_lane8_strm0 [0:4095];
  reg [31:0] pe37_lane8_strm0_tmp     ;
  reg [31:0] pe37_lane8_strm1 [0:4095];
  reg [31:0] pe37_lane8_strm1_tmp     ;
  reg [31:0] pe37_lane9_strm0 [0:4095];
  reg [31:0] pe37_lane9_strm0_tmp     ;
  reg [31:0] pe37_lane9_strm1 [0:4095];
  reg [31:0] pe37_lane9_strm1_tmp     ;
  reg [31:0] pe37_lane10_strm0 [0:4095];
  reg [31:0] pe37_lane10_strm0_tmp     ;
  reg [31:0] pe37_lane10_strm1 [0:4095];
  reg [31:0] pe37_lane10_strm1_tmp     ;
  reg [31:0] pe37_lane11_strm0 [0:4095];
  reg [31:0] pe37_lane11_strm0_tmp     ;
  reg [31:0] pe37_lane11_strm1 [0:4095];
  reg [31:0] pe37_lane11_strm1_tmp     ;
  reg [31:0] pe37_lane12_strm0 [0:4095];
  reg [31:0] pe37_lane12_strm0_tmp     ;
  reg [31:0] pe37_lane12_strm1 [0:4095];
  reg [31:0] pe37_lane12_strm1_tmp     ;
  reg [31:0] pe37_lane13_strm0 [0:4095];
  reg [31:0] pe37_lane13_strm0_tmp     ;
  reg [31:0] pe37_lane13_strm1 [0:4095];
  reg [31:0] pe37_lane13_strm1_tmp     ;
  reg [31:0] pe37_lane14_strm0 [0:4095];
  reg [31:0] pe37_lane14_strm0_tmp     ;
  reg [31:0] pe37_lane14_strm1 [0:4095];
  reg [31:0] pe37_lane14_strm1_tmp     ;
  reg [31:0] pe37_lane15_strm0 [0:4095];
  reg [31:0] pe37_lane15_strm0_tmp     ;
  reg [31:0] pe37_lane15_strm1 [0:4095];
  reg [31:0] pe37_lane15_strm1_tmp     ;
  reg [31:0] pe37_lane16_strm0 [0:4095];
  reg [31:0] pe37_lane16_strm0_tmp     ;
  reg [31:0] pe37_lane16_strm1 [0:4095];
  reg [31:0] pe37_lane16_strm1_tmp     ;
  reg [31:0] pe37_lane17_strm0 [0:4095];
  reg [31:0] pe37_lane17_strm0_tmp     ;
  reg [31:0] pe37_lane17_strm1 [0:4095];
  reg [31:0] pe37_lane17_strm1_tmp     ;
  reg [31:0] pe37_lane18_strm0 [0:4095];
  reg [31:0] pe37_lane18_strm0_tmp     ;
  reg [31:0] pe37_lane18_strm1 [0:4095];
  reg [31:0] pe37_lane18_strm1_tmp     ;
  reg [31:0] pe37_lane19_strm0 [0:4095];
  reg [31:0] pe37_lane19_strm0_tmp     ;
  reg [31:0] pe37_lane19_strm1 [0:4095];
  reg [31:0] pe37_lane19_strm1_tmp     ;
  reg [31:0] pe37_lane20_strm0 [0:4095];
  reg [31:0] pe37_lane20_strm0_tmp     ;
  reg [31:0] pe37_lane20_strm1 [0:4095];
  reg [31:0] pe37_lane20_strm1_tmp     ;
  reg [31:0] pe37_lane21_strm0 [0:4095];
  reg [31:0] pe37_lane21_strm0_tmp     ;
  reg [31:0] pe37_lane21_strm1 [0:4095];
  reg [31:0] pe37_lane21_strm1_tmp     ;
  reg [31:0] pe37_lane22_strm0 [0:4095];
  reg [31:0] pe37_lane22_strm0_tmp     ;
  reg [31:0] pe37_lane22_strm1 [0:4095];
  reg [31:0] pe37_lane22_strm1_tmp     ;
  reg [31:0] pe37_lane23_strm0 [0:4095];
  reg [31:0] pe37_lane23_strm0_tmp     ;
  reg [31:0] pe37_lane23_strm1 [0:4095];
  reg [31:0] pe37_lane23_strm1_tmp     ;
  reg [31:0] pe37_lane24_strm0 [0:4095];
  reg [31:0] pe37_lane24_strm0_tmp     ;
  reg [31:0] pe37_lane24_strm1 [0:4095];
  reg [31:0] pe37_lane24_strm1_tmp     ;
  reg [31:0] pe37_lane25_strm0 [0:4095];
  reg [31:0] pe37_lane25_strm0_tmp     ;
  reg [31:0] pe37_lane25_strm1 [0:4095];
  reg [31:0] pe37_lane25_strm1_tmp     ;
  reg [31:0] pe37_lane26_strm0 [0:4095];
  reg [31:0] pe37_lane26_strm0_tmp     ;
  reg [31:0] pe37_lane26_strm1 [0:4095];
  reg [31:0] pe37_lane26_strm1_tmp     ;
  reg [31:0] pe37_lane27_strm0 [0:4095];
  reg [31:0] pe37_lane27_strm0_tmp     ;
  reg [31:0] pe37_lane27_strm1 [0:4095];
  reg [31:0] pe37_lane27_strm1_tmp     ;
  reg [31:0] pe37_lane28_strm0 [0:4095];
  reg [31:0] pe37_lane28_strm0_tmp     ;
  reg [31:0] pe37_lane28_strm1 [0:4095];
  reg [31:0] pe37_lane28_strm1_tmp     ;
  reg [31:0] pe37_lane29_strm0 [0:4095];
  reg [31:0] pe37_lane29_strm0_tmp     ;
  reg [31:0] pe37_lane29_strm1 [0:4095];
  reg [31:0] pe37_lane29_strm1_tmp     ;
  reg [31:0] pe37_lane30_strm0 [0:4095];
  reg [31:0] pe37_lane30_strm0_tmp     ;
  reg [31:0] pe37_lane30_strm1 [0:4095];
  reg [31:0] pe37_lane30_strm1_tmp     ;
  reg [31:0] pe37_lane31_strm0 [0:4095];
  reg [31:0] pe37_lane31_strm0_tmp     ;
  reg [31:0] pe37_lane31_strm1 [0:4095];
  reg [31:0] pe37_lane31_strm1_tmp     ;
  reg [31:0] pe38_lane0_strm0 [0:4095];
  reg [31:0] pe38_lane0_strm0_tmp     ;
  reg [31:0] pe38_lane0_strm1 [0:4095];
  reg [31:0] pe38_lane0_strm1_tmp     ;
  reg [31:0] pe38_lane1_strm0 [0:4095];
  reg [31:0] pe38_lane1_strm0_tmp     ;
  reg [31:0] pe38_lane1_strm1 [0:4095];
  reg [31:0] pe38_lane1_strm1_tmp     ;
  reg [31:0] pe38_lane2_strm0 [0:4095];
  reg [31:0] pe38_lane2_strm0_tmp     ;
  reg [31:0] pe38_lane2_strm1 [0:4095];
  reg [31:0] pe38_lane2_strm1_tmp     ;
  reg [31:0] pe38_lane3_strm0 [0:4095];
  reg [31:0] pe38_lane3_strm0_tmp     ;
  reg [31:0] pe38_lane3_strm1 [0:4095];
  reg [31:0] pe38_lane3_strm1_tmp     ;
  reg [31:0] pe38_lane4_strm0 [0:4095];
  reg [31:0] pe38_lane4_strm0_tmp     ;
  reg [31:0] pe38_lane4_strm1 [0:4095];
  reg [31:0] pe38_lane4_strm1_tmp     ;
  reg [31:0] pe38_lane5_strm0 [0:4095];
  reg [31:0] pe38_lane5_strm0_tmp     ;
  reg [31:0] pe38_lane5_strm1 [0:4095];
  reg [31:0] pe38_lane5_strm1_tmp     ;
  reg [31:0] pe38_lane6_strm0 [0:4095];
  reg [31:0] pe38_lane6_strm0_tmp     ;
  reg [31:0] pe38_lane6_strm1 [0:4095];
  reg [31:0] pe38_lane6_strm1_tmp     ;
  reg [31:0] pe38_lane7_strm0 [0:4095];
  reg [31:0] pe38_lane7_strm0_tmp     ;
  reg [31:0] pe38_lane7_strm1 [0:4095];
  reg [31:0] pe38_lane7_strm1_tmp     ;
  reg [31:0] pe38_lane8_strm0 [0:4095];
  reg [31:0] pe38_lane8_strm0_tmp     ;
  reg [31:0] pe38_lane8_strm1 [0:4095];
  reg [31:0] pe38_lane8_strm1_tmp     ;
  reg [31:0] pe38_lane9_strm0 [0:4095];
  reg [31:0] pe38_lane9_strm0_tmp     ;
  reg [31:0] pe38_lane9_strm1 [0:4095];
  reg [31:0] pe38_lane9_strm1_tmp     ;
  reg [31:0] pe38_lane10_strm0 [0:4095];
  reg [31:0] pe38_lane10_strm0_tmp     ;
  reg [31:0] pe38_lane10_strm1 [0:4095];
  reg [31:0] pe38_lane10_strm1_tmp     ;
  reg [31:0] pe38_lane11_strm0 [0:4095];
  reg [31:0] pe38_lane11_strm0_tmp     ;
  reg [31:0] pe38_lane11_strm1 [0:4095];
  reg [31:0] pe38_lane11_strm1_tmp     ;
  reg [31:0] pe38_lane12_strm0 [0:4095];
  reg [31:0] pe38_lane12_strm0_tmp     ;
  reg [31:0] pe38_lane12_strm1 [0:4095];
  reg [31:0] pe38_lane12_strm1_tmp     ;
  reg [31:0] pe38_lane13_strm0 [0:4095];
  reg [31:0] pe38_lane13_strm0_tmp     ;
  reg [31:0] pe38_lane13_strm1 [0:4095];
  reg [31:0] pe38_lane13_strm1_tmp     ;
  reg [31:0] pe38_lane14_strm0 [0:4095];
  reg [31:0] pe38_lane14_strm0_tmp     ;
  reg [31:0] pe38_lane14_strm1 [0:4095];
  reg [31:0] pe38_lane14_strm1_tmp     ;
  reg [31:0] pe38_lane15_strm0 [0:4095];
  reg [31:0] pe38_lane15_strm0_tmp     ;
  reg [31:0] pe38_lane15_strm1 [0:4095];
  reg [31:0] pe38_lane15_strm1_tmp     ;
  reg [31:0] pe38_lane16_strm0 [0:4095];
  reg [31:0] pe38_lane16_strm0_tmp     ;
  reg [31:0] pe38_lane16_strm1 [0:4095];
  reg [31:0] pe38_lane16_strm1_tmp     ;
  reg [31:0] pe38_lane17_strm0 [0:4095];
  reg [31:0] pe38_lane17_strm0_tmp     ;
  reg [31:0] pe38_lane17_strm1 [0:4095];
  reg [31:0] pe38_lane17_strm1_tmp     ;
  reg [31:0] pe38_lane18_strm0 [0:4095];
  reg [31:0] pe38_lane18_strm0_tmp     ;
  reg [31:0] pe38_lane18_strm1 [0:4095];
  reg [31:0] pe38_lane18_strm1_tmp     ;
  reg [31:0] pe38_lane19_strm0 [0:4095];
  reg [31:0] pe38_lane19_strm0_tmp     ;
  reg [31:0] pe38_lane19_strm1 [0:4095];
  reg [31:0] pe38_lane19_strm1_tmp     ;
  reg [31:0] pe38_lane20_strm0 [0:4095];
  reg [31:0] pe38_lane20_strm0_tmp     ;
  reg [31:0] pe38_lane20_strm1 [0:4095];
  reg [31:0] pe38_lane20_strm1_tmp     ;
  reg [31:0] pe38_lane21_strm0 [0:4095];
  reg [31:0] pe38_lane21_strm0_tmp     ;
  reg [31:0] pe38_lane21_strm1 [0:4095];
  reg [31:0] pe38_lane21_strm1_tmp     ;
  reg [31:0] pe38_lane22_strm0 [0:4095];
  reg [31:0] pe38_lane22_strm0_tmp     ;
  reg [31:0] pe38_lane22_strm1 [0:4095];
  reg [31:0] pe38_lane22_strm1_tmp     ;
  reg [31:0] pe38_lane23_strm0 [0:4095];
  reg [31:0] pe38_lane23_strm0_tmp     ;
  reg [31:0] pe38_lane23_strm1 [0:4095];
  reg [31:0] pe38_lane23_strm1_tmp     ;
  reg [31:0] pe38_lane24_strm0 [0:4095];
  reg [31:0] pe38_lane24_strm0_tmp     ;
  reg [31:0] pe38_lane24_strm1 [0:4095];
  reg [31:0] pe38_lane24_strm1_tmp     ;
  reg [31:0] pe38_lane25_strm0 [0:4095];
  reg [31:0] pe38_lane25_strm0_tmp     ;
  reg [31:0] pe38_lane25_strm1 [0:4095];
  reg [31:0] pe38_lane25_strm1_tmp     ;
  reg [31:0] pe38_lane26_strm0 [0:4095];
  reg [31:0] pe38_lane26_strm0_tmp     ;
  reg [31:0] pe38_lane26_strm1 [0:4095];
  reg [31:0] pe38_lane26_strm1_tmp     ;
  reg [31:0] pe38_lane27_strm0 [0:4095];
  reg [31:0] pe38_lane27_strm0_tmp     ;
  reg [31:0] pe38_lane27_strm1 [0:4095];
  reg [31:0] pe38_lane27_strm1_tmp     ;
  reg [31:0] pe38_lane28_strm0 [0:4095];
  reg [31:0] pe38_lane28_strm0_tmp     ;
  reg [31:0] pe38_lane28_strm1 [0:4095];
  reg [31:0] pe38_lane28_strm1_tmp     ;
  reg [31:0] pe38_lane29_strm0 [0:4095];
  reg [31:0] pe38_lane29_strm0_tmp     ;
  reg [31:0] pe38_lane29_strm1 [0:4095];
  reg [31:0] pe38_lane29_strm1_tmp     ;
  reg [31:0] pe38_lane30_strm0 [0:4095];
  reg [31:0] pe38_lane30_strm0_tmp     ;
  reg [31:0] pe38_lane30_strm1 [0:4095];
  reg [31:0] pe38_lane30_strm1_tmp     ;
  reg [31:0] pe38_lane31_strm0 [0:4095];
  reg [31:0] pe38_lane31_strm0_tmp     ;
  reg [31:0] pe38_lane31_strm1 [0:4095];
  reg [31:0] pe38_lane31_strm1_tmp     ;
  reg [31:0] pe39_lane0_strm0 [0:4095];
  reg [31:0] pe39_lane0_strm0_tmp     ;
  reg [31:0] pe39_lane0_strm1 [0:4095];
  reg [31:0] pe39_lane0_strm1_tmp     ;
  reg [31:0] pe39_lane1_strm0 [0:4095];
  reg [31:0] pe39_lane1_strm0_tmp     ;
  reg [31:0] pe39_lane1_strm1 [0:4095];
  reg [31:0] pe39_lane1_strm1_tmp     ;
  reg [31:0] pe39_lane2_strm0 [0:4095];
  reg [31:0] pe39_lane2_strm0_tmp     ;
  reg [31:0] pe39_lane2_strm1 [0:4095];
  reg [31:0] pe39_lane2_strm1_tmp     ;
  reg [31:0] pe39_lane3_strm0 [0:4095];
  reg [31:0] pe39_lane3_strm0_tmp     ;
  reg [31:0] pe39_lane3_strm1 [0:4095];
  reg [31:0] pe39_lane3_strm1_tmp     ;
  reg [31:0] pe39_lane4_strm0 [0:4095];
  reg [31:0] pe39_lane4_strm0_tmp     ;
  reg [31:0] pe39_lane4_strm1 [0:4095];
  reg [31:0] pe39_lane4_strm1_tmp     ;
  reg [31:0] pe39_lane5_strm0 [0:4095];
  reg [31:0] pe39_lane5_strm0_tmp     ;
  reg [31:0] pe39_lane5_strm1 [0:4095];
  reg [31:0] pe39_lane5_strm1_tmp     ;
  reg [31:0] pe39_lane6_strm0 [0:4095];
  reg [31:0] pe39_lane6_strm0_tmp     ;
  reg [31:0] pe39_lane6_strm1 [0:4095];
  reg [31:0] pe39_lane6_strm1_tmp     ;
  reg [31:0] pe39_lane7_strm0 [0:4095];
  reg [31:0] pe39_lane7_strm0_tmp     ;
  reg [31:0] pe39_lane7_strm1 [0:4095];
  reg [31:0] pe39_lane7_strm1_tmp     ;
  reg [31:0] pe39_lane8_strm0 [0:4095];
  reg [31:0] pe39_lane8_strm0_tmp     ;
  reg [31:0] pe39_lane8_strm1 [0:4095];
  reg [31:0] pe39_lane8_strm1_tmp     ;
  reg [31:0] pe39_lane9_strm0 [0:4095];
  reg [31:0] pe39_lane9_strm0_tmp     ;
  reg [31:0] pe39_lane9_strm1 [0:4095];
  reg [31:0] pe39_lane9_strm1_tmp     ;
  reg [31:0] pe39_lane10_strm0 [0:4095];
  reg [31:0] pe39_lane10_strm0_tmp     ;
  reg [31:0] pe39_lane10_strm1 [0:4095];
  reg [31:0] pe39_lane10_strm1_tmp     ;
  reg [31:0] pe39_lane11_strm0 [0:4095];
  reg [31:0] pe39_lane11_strm0_tmp     ;
  reg [31:0] pe39_lane11_strm1 [0:4095];
  reg [31:0] pe39_lane11_strm1_tmp     ;
  reg [31:0] pe39_lane12_strm0 [0:4095];
  reg [31:0] pe39_lane12_strm0_tmp     ;
  reg [31:0] pe39_lane12_strm1 [0:4095];
  reg [31:0] pe39_lane12_strm1_tmp     ;
  reg [31:0] pe39_lane13_strm0 [0:4095];
  reg [31:0] pe39_lane13_strm0_tmp     ;
  reg [31:0] pe39_lane13_strm1 [0:4095];
  reg [31:0] pe39_lane13_strm1_tmp     ;
  reg [31:0] pe39_lane14_strm0 [0:4095];
  reg [31:0] pe39_lane14_strm0_tmp     ;
  reg [31:0] pe39_lane14_strm1 [0:4095];
  reg [31:0] pe39_lane14_strm1_tmp     ;
  reg [31:0] pe39_lane15_strm0 [0:4095];
  reg [31:0] pe39_lane15_strm0_tmp     ;
  reg [31:0] pe39_lane15_strm1 [0:4095];
  reg [31:0] pe39_lane15_strm1_tmp     ;
  reg [31:0] pe39_lane16_strm0 [0:4095];
  reg [31:0] pe39_lane16_strm0_tmp     ;
  reg [31:0] pe39_lane16_strm1 [0:4095];
  reg [31:0] pe39_lane16_strm1_tmp     ;
  reg [31:0] pe39_lane17_strm0 [0:4095];
  reg [31:0] pe39_lane17_strm0_tmp     ;
  reg [31:0] pe39_lane17_strm1 [0:4095];
  reg [31:0] pe39_lane17_strm1_tmp     ;
  reg [31:0] pe39_lane18_strm0 [0:4095];
  reg [31:0] pe39_lane18_strm0_tmp     ;
  reg [31:0] pe39_lane18_strm1 [0:4095];
  reg [31:0] pe39_lane18_strm1_tmp     ;
  reg [31:0] pe39_lane19_strm0 [0:4095];
  reg [31:0] pe39_lane19_strm0_tmp     ;
  reg [31:0] pe39_lane19_strm1 [0:4095];
  reg [31:0] pe39_lane19_strm1_tmp     ;
  reg [31:0] pe39_lane20_strm0 [0:4095];
  reg [31:0] pe39_lane20_strm0_tmp     ;
  reg [31:0] pe39_lane20_strm1 [0:4095];
  reg [31:0] pe39_lane20_strm1_tmp     ;
  reg [31:0] pe39_lane21_strm0 [0:4095];
  reg [31:0] pe39_lane21_strm0_tmp     ;
  reg [31:0] pe39_lane21_strm1 [0:4095];
  reg [31:0] pe39_lane21_strm1_tmp     ;
  reg [31:0] pe39_lane22_strm0 [0:4095];
  reg [31:0] pe39_lane22_strm0_tmp     ;
  reg [31:0] pe39_lane22_strm1 [0:4095];
  reg [31:0] pe39_lane22_strm1_tmp     ;
  reg [31:0] pe39_lane23_strm0 [0:4095];
  reg [31:0] pe39_lane23_strm0_tmp     ;
  reg [31:0] pe39_lane23_strm1 [0:4095];
  reg [31:0] pe39_lane23_strm1_tmp     ;
  reg [31:0] pe39_lane24_strm0 [0:4095];
  reg [31:0] pe39_lane24_strm0_tmp     ;
  reg [31:0] pe39_lane24_strm1 [0:4095];
  reg [31:0] pe39_lane24_strm1_tmp     ;
  reg [31:0] pe39_lane25_strm0 [0:4095];
  reg [31:0] pe39_lane25_strm0_tmp     ;
  reg [31:0] pe39_lane25_strm1 [0:4095];
  reg [31:0] pe39_lane25_strm1_tmp     ;
  reg [31:0] pe39_lane26_strm0 [0:4095];
  reg [31:0] pe39_lane26_strm0_tmp     ;
  reg [31:0] pe39_lane26_strm1 [0:4095];
  reg [31:0] pe39_lane26_strm1_tmp     ;
  reg [31:0] pe39_lane27_strm0 [0:4095];
  reg [31:0] pe39_lane27_strm0_tmp     ;
  reg [31:0] pe39_lane27_strm1 [0:4095];
  reg [31:0] pe39_lane27_strm1_tmp     ;
  reg [31:0] pe39_lane28_strm0 [0:4095];
  reg [31:0] pe39_lane28_strm0_tmp     ;
  reg [31:0] pe39_lane28_strm1 [0:4095];
  reg [31:0] pe39_lane28_strm1_tmp     ;
  reg [31:0] pe39_lane29_strm0 [0:4095];
  reg [31:0] pe39_lane29_strm0_tmp     ;
  reg [31:0] pe39_lane29_strm1 [0:4095];
  reg [31:0] pe39_lane29_strm1_tmp     ;
  reg [31:0] pe39_lane30_strm0 [0:4095];
  reg [31:0] pe39_lane30_strm0_tmp     ;
  reg [31:0] pe39_lane30_strm1 [0:4095];
  reg [31:0] pe39_lane30_strm1_tmp     ;
  reg [31:0] pe39_lane31_strm0 [0:4095];
  reg [31:0] pe39_lane31_strm0_tmp     ;
  reg [31:0] pe39_lane31_strm1 [0:4095];
  reg [31:0] pe39_lane31_strm1_tmp     ;
  reg [31:0] pe40_lane0_strm0 [0:4095];
  reg [31:0] pe40_lane0_strm0_tmp     ;
  reg [31:0] pe40_lane0_strm1 [0:4095];
  reg [31:0] pe40_lane0_strm1_tmp     ;
  reg [31:0] pe40_lane1_strm0 [0:4095];
  reg [31:0] pe40_lane1_strm0_tmp     ;
  reg [31:0] pe40_lane1_strm1 [0:4095];
  reg [31:0] pe40_lane1_strm1_tmp     ;
  reg [31:0] pe40_lane2_strm0 [0:4095];
  reg [31:0] pe40_lane2_strm0_tmp     ;
  reg [31:0] pe40_lane2_strm1 [0:4095];
  reg [31:0] pe40_lane2_strm1_tmp     ;
  reg [31:0] pe40_lane3_strm0 [0:4095];
  reg [31:0] pe40_lane3_strm0_tmp     ;
  reg [31:0] pe40_lane3_strm1 [0:4095];
  reg [31:0] pe40_lane3_strm1_tmp     ;
  reg [31:0] pe40_lane4_strm0 [0:4095];
  reg [31:0] pe40_lane4_strm0_tmp     ;
  reg [31:0] pe40_lane4_strm1 [0:4095];
  reg [31:0] pe40_lane4_strm1_tmp     ;
  reg [31:0] pe40_lane5_strm0 [0:4095];
  reg [31:0] pe40_lane5_strm0_tmp     ;
  reg [31:0] pe40_lane5_strm1 [0:4095];
  reg [31:0] pe40_lane5_strm1_tmp     ;
  reg [31:0] pe40_lane6_strm0 [0:4095];
  reg [31:0] pe40_lane6_strm0_tmp     ;
  reg [31:0] pe40_lane6_strm1 [0:4095];
  reg [31:0] pe40_lane6_strm1_tmp     ;
  reg [31:0] pe40_lane7_strm0 [0:4095];
  reg [31:0] pe40_lane7_strm0_tmp     ;
  reg [31:0] pe40_lane7_strm1 [0:4095];
  reg [31:0] pe40_lane7_strm1_tmp     ;
  reg [31:0] pe40_lane8_strm0 [0:4095];
  reg [31:0] pe40_lane8_strm0_tmp     ;
  reg [31:0] pe40_lane8_strm1 [0:4095];
  reg [31:0] pe40_lane8_strm1_tmp     ;
  reg [31:0] pe40_lane9_strm0 [0:4095];
  reg [31:0] pe40_lane9_strm0_tmp     ;
  reg [31:0] pe40_lane9_strm1 [0:4095];
  reg [31:0] pe40_lane9_strm1_tmp     ;
  reg [31:0] pe40_lane10_strm0 [0:4095];
  reg [31:0] pe40_lane10_strm0_tmp     ;
  reg [31:0] pe40_lane10_strm1 [0:4095];
  reg [31:0] pe40_lane10_strm1_tmp     ;
  reg [31:0] pe40_lane11_strm0 [0:4095];
  reg [31:0] pe40_lane11_strm0_tmp     ;
  reg [31:0] pe40_lane11_strm1 [0:4095];
  reg [31:0] pe40_lane11_strm1_tmp     ;
  reg [31:0] pe40_lane12_strm0 [0:4095];
  reg [31:0] pe40_lane12_strm0_tmp     ;
  reg [31:0] pe40_lane12_strm1 [0:4095];
  reg [31:0] pe40_lane12_strm1_tmp     ;
  reg [31:0] pe40_lane13_strm0 [0:4095];
  reg [31:0] pe40_lane13_strm0_tmp     ;
  reg [31:0] pe40_lane13_strm1 [0:4095];
  reg [31:0] pe40_lane13_strm1_tmp     ;
  reg [31:0] pe40_lane14_strm0 [0:4095];
  reg [31:0] pe40_lane14_strm0_tmp     ;
  reg [31:0] pe40_lane14_strm1 [0:4095];
  reg [31:0] pe40_lane14_strm1_tmp     ;
  reg [31:0] pe40_lane15_strm0 [0:4095];
  reg [31:0] pe40_lane15_strm0_tmp     ;
  reg [31:0] pe40_lane15_strm1 [0:4095];
  reg [31:0] pe40_lane15_strm1_tmp     ;
  reg [31:0] pe40_lane16_strm0 [0:4095];
  reg [31:0] pe40_lane16_strm0_tmp     ;
  reg [31:0] pe40_lane16_strm1 [0:4095];
  reg [31:0] pe40_lane16_strm1_tmp     ;
  reg [31:0] pe40_lane17_strm0 [0:4095];
  reg [31:0] pe40_lane17_strm0_tmp     ;
  reg [31:0] pe40_lane17_strm1 [0:4095];
  reg [31:0] pe40_lane17_strm1_tmp     ;
  reg [31:0] pe40_lane18_strm0 [0:4095];
  reg [31:0] pe40_lane18_strm0_tmp     ;
  reg [31:0] pe40_lane18_strm1 [0:4095];
  reg [31:0] pe40_lane18_strm1_tmp     ;
  reg [31:0] pe40_lane19_strm0 [0:4095];
  reg [31:0] pe40_lane19_strm0_tmp     ;
  reg [31:0] pe40_lane19_strm1 [0:4095];
  reg [31:0] pe40_lane19_strm1_tmp     ;
  reg [31:0] pe40_lane20_strm0 [0:4095];
  reg [31:0] pe40_lane20_strm0_tmp     ;
  reg [31:0] pe40_lane20_strm1 [0:4095];
  reg [31:0] pe40_lane20_strm1_tmp     ;
  reg [31:0] pe40_lane21_strm0 [0:4095];
  reg [31:0] pe40_lane21_strm0_tmp     ;
  reg [31:0] pe40_lane21_strm1 [0:4095];
  reg [31:0] pe40_lane21_strm1_tmp     ;
  reg [31:0] pe40_lane22_strm0 [0:4095];
  reg [31:0] pe40_lane22_strm0_tmp     ;
  reg [31:0] pe40_lane22_strm1 [0:4095];
  reg [31:0] pe40_lane22_strm1_tmp     ;
  reg [31:0] pe40_lane23_strm0 [0:4095];
  reg [31:0] pe40_lane23_strm0_tmp     ;
  reg [31:0] pe40_lane23_strm1 [0:4095];
  reg [31:0] pe40_lane23_strm1_tmp     ;
  reg [31:0] pe40_lane24_strm0 [0:4095];
  reg [31:0] pe40_lane24_strm0_tmp     ;
  reg [31:0] pe40_lane24_strm1 [0:4095];
  reg [31:0] pe40_lane24_strm1_tmp     ;
  reg [31:0] pe40_lane25_strm0 [0:4095];
  reg [31:0] pe40_lane25_strm0_tmp     ;
  reg [31:0] pe40_lane25_strm1 [0:4095];
  reg [31:0] pe40_lane25_strm1_tmp     ;
  reg [31:0] pe40_lane26_strm0 [0:4095];
  reg [31:0] pe40_lane26_strm0_tmp     ;
  reg [31:0] pe40_lane26_strm1 [0:4095];
  reg [31:0] pe40_lane26_strm1_tmp     ;
  reg [31:0] pe40_lane27_strm0 [0:4095];
  reg [31:0] pe40_lane27_strm0_tmp     ;
  reg [31:0] pe40_lane27_strm1 [0:4095];
  reg [31:0] pe40_lane27_strm1_tmp     ;
  reg [31:0] pe40_lane28_strm0 [0:4095];
  reg [31:0] pe40_lane28_strm0_tmp     ;
  reg [31:0] pe40_lane28_strm1 [0:4095];
  reg [31:0] pe40_lane28_strm1_tmp     ;
  reg [31:0] pe40_lane29_strm0 [0:4095];
  reg [31:0] pe40_lane29_strm0_tmp     ;
  reg [31:0] pe40_lane29_strm1 [0:4095];
  reg [31:0] pe40_lane29_strm1_tmp     ;
  reg [31:0] pe40_lane30_strm0 [0:4095];
  reg [31:0] pe40_lane30_strm0_tmp     ;
  reg [31:0] pe40_lane30_strm1 [0:4095];
  reg [31:0] pe40_lane30_strm1_tmp     ;
  reg [31:0] pe40_lane31_strm0 [0:4095];
  reg [31:0] pe40_lane31_strm0_tmp     ;
  reg [31:0] pe40_lane31_strm1 [0:4095];
  reg [31:0] pe40_lane31_strm1_tmp     ;
  reg [31:0] pe41_lane0_strm0 [0:4095];
  reg [31:0] pe41_lane0_strm0_tmp     ;
  reg [31:0] pe41_lane0_strm1 [0:4095];
  reg [31:0] pe41_lane0_strm1_tmp     ;
  reg [31:0] pe41_lane1_strm0 [0:4095];
  reg [31:0] pe41_lane1_strm0_tmp     ;
  reg [31:0] pe41_lane1_strm1 [0:4095];
  reg [31:0] pe41_lane1_strm1_tmp     ;
  reg [31:0] pe41_lane2_strm0 [0:4095];
  reg [31:0] pe41_lane2_strm0_tmp     ;
  reg [31:0] pe41_lane2_strm1 [0:4095];
  reg [31:0] pe41_lane2_strm1_tmp     ;
  reg [31:0] pe41_lane3_strm0 [0:4095];
  reg [31:0] pe41_lane3_strm0_tmp     ;
  reg [31:0] pe41_lane3_strm1 [0:4095];
  reg [31:0] pe41_lane3_strm1_tmp     ;
  reg [31:0] pe41_lane4_strm0 [0:4095];
  reg [31:0] pe41_lane4_strm0_tmp     ;
  reg [31:0] pe41_lane4_strm1 [0:4095];
  reg [31:0] pe41_lane4_strm1_tmp     ;
  reg [31:0] pe41_lane5_strm0 [0:4095];
  reg [31:0] pe41_lane5_strm0_tmp     ;
  reg [31:0] pe41_lane5_strm1 [0:4095];
  reg [31:0] pe41_lane5_strm1_tmp     ;
  reg [31:0] pe41_lane6_strm0 [0:4095];
  reg [31:0] pe41_lane6_strm0_tmp     ;
  reg [31:0] pe41_lane6_strm1 [0:4095];
  reg [31:0] pe41_lane6_strm1_tmp     ;
  reg [31:0] pe41_lane7_strm0 [0:4095];
  reg [31:0] pe41_lane7_strm0_tmp     ;
  reg [31:0] pe41_lane7_strm1 [0:4095];
  reg [31:0] pe41_lane7_strm1_tmp     ;
  reg [31:0] pe41_lane8_strm0 [0:4095];
  reg [31:0] pe41_lane8_strm0_tmp     ;
  reg [31:0] pe41_lane8_strm1 [0:4095];
  reg [31:0] pe41_lane8_strm1_tmp     ;
  reg [31:0] pe41_lane9_strm0 [0:4095];
  reg [31:0] pe41_lane9_strm0_tmp     ;
  reg [31:0] pe41_lane9_strm1 [0:4095];
  reg [31:0] pe41_lane9_strm1_tmp     ;
  reg [31:0] pe41_lane10_strm0 [0:4095];
  reg [31:0] pe41_lane10_strm0_tmp     ;
  reg [31:0] pe41_lane10_strm1 [0:4095];
  reg [31:0] pe41_lane10_strm1_tmp     ;
  reg [31:0] pe41_lane11_strm0 [0:4095];
  reg [31:0] pe41_lane11_strm0_tmp     ;
  reg [31:0] pe41_lane11_strm1 [0:4095];
  reg [31:0] pe41_lane11_strm1_tmp     ;
  reg [31:0] pe41_lane12_strm0 [0:4095];
  reg [31:0] pe41_lane12_strm0_tmp     ;
  reg [31:0] pe41_lane12_strm1 [0:4095];
  reg [31:0] pe41_lane12_strm1_tmp     ;
  reg [31:0] pe41_lane13_strm0 [0:4095];
  reg [31:0] pe41_lane13_strm0_tmp     ;
  reg [31:0] pe41_lane13_strm1 [0:4095];
  reg [31:0] pe41_lane13_strm1_tmp     ;
  reg [31:0] pe41_lane14_strm0 [0:4095];
  reg [31:0] pe41_lane14_strm0_tmp     ;
  reg [31:0] pe41_lane14_strm1 [0:4095];
  reg [31:0] pe41_lane14_strm1_tmp     ;
  reg [31:0] pe41_lane15_strm0 [0:4095];
  reg [31:0] pe41_lane15_strm0_tmp     ;
  reg [31:0] pe41_lane15_strm1 [0:4095];
  reg [31:0] pe41_lane15_strm1_tmp     ;
  reg [31:0] pe41_lane16_strm0 [0:4095];
  reg [31:0] pe41_lane16_strm0_tmp     ;
  reg [31:0] pe41_lane16_strm1 [0:4095];
  reg [31:0] pe41_lane16_strm1_tmp     ;
  reg [31:0] pe41_lane17_strm0 [0:4095];
  reg [31:0] pe41_lane17_strm0_tmp     ;
  reg [31:0] pe41_lane17_strm1 [0:4095];
  reg [31:0] pe41_lane17_strm1_tmp     ;
  reg [31:0] pe41_lane18_strm0 [0:4095];
  reg [31:0] pe41_lane18_strm0_tmp     ;
  reg [31:0] pe41_lane18_strm1 [0:4095];
  reg [31:0] pe41_lane18_strm1_tmp     ;
  reg [31:0] pe41_lane19_strm0 [0:4095];
  reg [31:0] pe41_lane19_strm0_tmp     ;
  reg [31:0] pe41_lane19_strm1 [0:4095];
  reg [31:0] pe41_lane19_strm1_tmp     ;
  reg [31:0] pe41_lane20_strm0 [0:4095];
  reg [31:0] pe41_lane20_strm0_tmp     ;
  reg [31:0] pe41_lane20_strm1 [0:4095];
  reg [31:0] pe41_lane20_strm1_tmp     ;
  reg [31:0] pe41_lane21_strm0 [0:4095];
  reg [31:0] pe41_lane21_strm0_tmp     ;
  reg [31:0] pe41_lane21_strm1 [0:4095];
  reg [31:0] pe41_lane21_strm1_tmp     ;
  reg [31:0] pe41_lane22_strm0 [0:4095];
  reg [31:0] pe41_lane22_strm0_tmp     ;
  reg [31:0] pe41_lane22_strm1 [0:4095];
  reg [31:0] pe41_lane22_strm1_tmp     ;
  reg [31:0] pe41_lane23_strm0 [0:4095];
  reg [31:0] pe41_lane23_strm0_tmp     ;
  reg [31:0] pe41_lane23_strm1 [0:4095];
  reg [31:0] pe41_lane23_strm1_tmp     ;
  reg [31:0] pe41_lane24_strm0 [0:4095];
  reg [31:0] pe41_lane24_strm0_tmp     ;
  reg [31:0] pe41_lane24_strm1 [0:4095];
  reg [31:0] pe41_lane24_strm1_tmp     ;
  reg [31:0] pe41_lane25_strm0 [0:4095];
  reg [31:0] pe41_lane25_strm0_tmp     ;
  reg [31:0] pe41_lane25_strm1 [0:4095];
  reg [31:0] pe41_lane25_strm1_tmp     ;
  reg [31:0] pe41_lane26_strm0 [0:4095];
  reg [31:0] pe41_lane26_strm0_tmp     ;
  reg [31:0] pe41_lane26_strm1 [0:4095];
  reg [31:0] pe41_lane26_strm1_tmp     ;
  reg [31:0] pe41_lane27_strm0 [0:4095];
  reg [31:0] pe41_lane27_strm0_tmp     ;
  reg [31:0] pe41_lane27_strm1 [0:4095];
  reg [31:0] pe41_lane27_strm1_tmp     ;
  reg [31:0] pe41_lane28_strm0 [0:4095];
  reg [31:0] pe41_lane28_strm0_tmp     ;
  reg [31:0] pe41_lane28_strm1 [0:4095];
  reg [31:0] pe41_lane28_strm1_tmp     ;
  reg [31:0] pe41_lane29_strm0 [0:4095];
  reg [31:0] pe41_lane29_strm0_tmp     ;
  reg [31:0] pe41_lane29_strm1 [0:4095];
  reg [31:0] pe41_lane29_strm1_tmp     ;
  reg [31:0] pe41_lane30_strm0 [0:4095];
  reg [31:0] pe41_lane30_strm0_tmp     ;
  reg [31:0] pe41_lane30_strm1 [0:4095];
  reg [31:0] pe41_lane30_strm1_tmp     ;
  reg [31:0] pe41_lane31_strm0 [0:4095];
  reg [31:0] pe41_lane31_strm0_tmp     ;
  reg [31:0] pe41_lane31_strm1 [0:4095];
  reg [31:0] pe41_lane31_strm1_tmp     ;
  reg [31:0] pe42_lane0_strm0 [0:4095];
  reg [31:0] pe42_lane0_strm0_tmp     ;
  reg [31:0] pe42_lane0_strm1 [0:4095];
  reg [31:0] pe42_lane0_strm1_tmp     ;
  reg [31:0] pe42_lane1_strm0 [0:4095];
  reg [31:0] pe42_lane1_strm0_tmp     ;
  reg [31:0] pe42_lane1_strm1 [0:4095];
  reg [31:0] pe42_lane1_strm1_tmp     ;
  reg [31:0] pe42_lane2_strm0 [0:4095];
  reg [31:0] pe42_lane2_strm0_tmp     ;
  reg [31:0] pe42_lane2_strm1 [0:4095];
  reg [31:0] pe42_lane2_strm1_tmp     ;
  reg [31:0] pe42_lane3_strm0 [0:4095];
  reg [31:0] pe42_lane3_strm0_tmp     ;
  reg [31:0] pe42_lane3_strm1 [0:4095];
  reg [31:0] pe42_lane3_strm1_tmp     ;
  reg [31:0] pe42_lane4_strm0 [0:4095];
  reg [31:0] pe42_lane4_strm0_tmp     ;
  reg [31:0] pe42_lane4_strm1 [0:4095];
  reg [31:0] pe42_lane4_strm1_tmp     ;
  reg [31:0] pe42_lane5_strm0 [0:4095];
  reg [31:0] pe42_lane5_strm0_tmp     ;
  reg [31:0] pe42_lane5_strm1 [0:4095];
  reg [31:0] pe42_lane5_strm1_tmp     ;
  reg [31:0] pe42_lane6_strm0 [0:4095];
  reg [31:0] pe42_lane6_strm0_tmp     ;
  reg [31:0] pe42_lane6_strm1 [0:4095];
  reg [31:0] pe42_lane6_strm1_tmp     ;
  reg [31:0] pe42_lane7_strm0 [0:4095];
  reg [31:0] pe42_lane7_strm0_tmp     ;
  reg [31:0] pe42_lane7_strm1 [0:4095];
  reg [31:0] pe42_lane7_strm1_tmp     ;
  reg [31:0] pe42_lane8_strm0 [0:4095];
  reg [31:0] pe42_lane8_strm0_tmp     ;
  reg [31:0] pe42_lane8_strm1 [0:4095];
  reg [31:0] pe42_lane8_strm1_tmp     ;
  reg [31:0] pe42_lane9_strm0 [0:4095];
  reg [31:0] pe42_lane9_strm0_tmp     ;
  reg [31:0] pe42_lane9_strm1 [0:4095];
  reg [31:0] pe42_lane9_strm1_tmp     ;
  reg [31:0] pe42_lane10_strm0 [0:4095];
  reg [31:0] pe42_lane10_strm0_tmp     ;
  reg [31:0] pe42_lane10_strm1 [0:4095];
  reg [31:0] pe42_lane10_strm1_tmp     ;
  reg [31:0] pe42_lane11_strm0 [0:4095];
  reg [31:0] pe42_lane11_strm0_tmp     ;
  reg [31:0] pe42_lane11_strm1 [0:4095];
  reg [31:0] pe42_lane11_strm1_tmp     ;
  reg [31:0] pe42_lane12_strm0 [0:4095];
  reg [31:0] pe42_lane12_strm0_tmp     ;
  reg [31:0] pe42_lane12_strm1 [0:4095];
  reg [31:0] pe42_lane12_strm1_tmp     ;
  reg [31:0] pe42_lane13_strm0 [0:4095];
  reg [31:0] pe42_lane13_strm0_tmp     ;
  reg [31:0] pe42_lane13_strm1 [0:4095];
  reg [31:0] pe42_lane13_strm1_tmp     ;
  reg [31:0] pe42_lane14_strm0 [0:4095];
  reg [31:0] pe42_lane14_strm0_tmp     ;
  reg [31:0] pe42_lane14_strm1 [0:4095];
  reg [31:0] pe42_lane14_strm1_tmp     ;
  reg [31:0] pe42_lane15_strm0 [0:4095];
  reg [31:0] pe42_lane15_strm0_tmp     ;
  reg [31:0] pe42_lane15_strm1 [0:4095];
  reg [31:0] pe42_lane15_strm1_tmp     ;
  reg [31:0] pe42_lane16_strm0 [0:4095];
  reg [31:0] pe42_lane16_strm0_tmp     ;
  reg [31:0] pe42_lane16_strm1 [0:4095];
  reg [31:0] pe42_lane16_strm1_tmp     ;
  reg [31:0] pe42_lane17_strm0 [0:4095];
  reg [31:0] pe42_lane17_strm0_tmp     ;
  reg [31:0] pe42_lane17_strm1 [0:4095];
  reg [31:0] pe42_lane17_strm1_tmp     ;
  reg [31:0] pe42_lane18_strm0 [0:4095];
  reg [31:0] pe42_lane18_strm0_tmp     ;
  reg [31:0] pe42_lane18_strm1 [0:4095];
  reg [31:0] pe42_lane18_strm1_tmp     ;
  reg [31:0] pe42_lane19_strm0 [0:4095];
  reg [31:0] pe42_lane19_strm0_tmp     ;
  reg [31:0] pe42_lane19_strm1 [0:4095];
  reg [31:0] pe42_lane19_strm1_tmp     ;
  reg [31:0] pe42_lane20_strm0 [0:4095];
  reg [31:0] pe42_lane20_strm0_tmp     ;
  reg [31:0] pe42_lane20_strm1 [0:4095];
  reg [31:0] pe42_lane20_strm1_tmp     ;
  reg [31:0] pe42_lane21_strm0 [0:4095];
  reg [31:0] pe42_lane21_strm0_tmp     ;
  reg [31:0] pe42_lane21_strm1 [0:4095];
  reg [31:0] pe42_lane21_strm1_tmp     ;
  reg [31:0] pe42_lane22_strm0 [0:4095];
  reg [31:0] pe42_lane22_strm0_tmp     ;
  reg [31:0] pe42_lane22_strm1 [0:4095];
  reg [31:0] pe42_lane22_strm1_tmp     ;
  reg [31:0] pe42_lane23_strm0 [0:4095];
  reg [31:0] pe42_lane23_strm0_tmp     ;
  reg [31:0] pe42_lane23_strm1 [0:4095];
  reg [31:0] pe42_lane23_strm1_tmp     ;
  reg [31:0] pe42_lane24_strm0 [0:4095];
  reg [31:0] pe42_lane24_strm0_tmp     ;
  reg [31:0] pe42_lane24_strm1 [0:4095];
  reg [31:0] pe42_lane24_strm1_tmp     ;
  reg [31:0] pe42_lane25_strm0 [0:4095];
  reg [31:0] pe42_lane25_strm0_tmp     ;
  reg [31:0] pe42_lane25_strm1 [0:4095];
  reg [31:0] pe42_lane25_strm1_tmp     ;
  reg [31:0] pe42_lane26_strm0 [0:4095];
  reg [31:0] pe42_lane26_strm0_tmp     ;
  reg [31:0] pe42_lane26_strm1 [0:4095];
  reg [31:0] pe42_lane26_strm1_tmp     ;
  reg [31:0] pe42_lane27_strm0 [0:4095];
  reg [31:0] pe42_lane27_strm0_tmp     ;
  reg [31:0] pe42_lane27_strm1 [0:4095];
  reg [31:0] pe42_lane27_strm1_tmp     ;
  reg [31:0] pe42_lane28_strm0 [0:4095];
  reg [31:0] pe42_lane28_strm0_tmp     ;
  reg [31:0] pe42_lane28_strm1 [0:4095];
  reg [31:0] pe42_lane28_strm1_tmp     ;
  reg [31:0] pe42_lane29_strm0 [0:4095];
  reg [31:0] pe42_lane29_strm0_tmp     ;
  reg [31:0] pe42_lane29_strm1 [0:4095];
  reg [31:0] pe42_lane29_strm1_tmp     ;
  reg [31:0] pe42_lane30_strm0 [0:4095];
  reg [31:0] pe42_lane30_strm0_tmp     ;
  reg [31:0] pe42_lane30_strm1 [0:4095];
  reg [31:0] pe42_lane30_strm1_tmp     ;
  reg [31:0] pe42_lane31_strm0 [0:4095];
  reg [31:0] pe42_lane31_strm0_tmp     ;
  reg [31:0] pe42_lane31_strm1 [0:4095];
  reg [31:0] pe42_lane31_strm1_tmp     ;
  reg [31:0] pe43_lane0_strm0 [0:4095];
  reg [31:0] pe43_lane0_strm0_tmp     ;
  reg [31:0] pe43_lane0_strm1 [0:4095];
  reg [31:0] pe43_lane0_strm1_tmp     ;
  reg [31:0] pe43_lane1_strm0 [0:4095];
  reg [31:0] pe43_lane1_strm0_tmp     ;
  reg [31:0] pe43_lane1_strm1 [0:4095];
  reg [31:0] pe43_lane1_strm1_tmp     ;
  reg [31:0] pe43_lane2_strm0 [0:4095];
  reg [31:0] pe43_lane2_strm0_tmp     ;
  reg [31:0] pe43_lane2_strm1 [0:4095];
  reg [31:0] pe43_lane2_strm1_tmp     ;
  reg [31:0] pe43_lane3_strm0 [0:4095];
  reg [31:0] pe43_lane3_strm0_tmp     ;
  reg [31:0] pe43_lane3_strm1 [0:4095];
  reg [31:0] pe43_lane3_strm1_tmp     ;
  reg [31:0] pe43_lane4_strm0 [0:4095];
  reg [31:0] pe43_lane4_strm0_tmp     ;
  reg [31:0] pe43_lane4_strm1 [0:4095];
  reg [31:0] pe43_lane4_strm1_tmp     ;
  reg [31:0] pe43_lane5_strm0 [0:4095];
  reg [31:0] pe43_lane5_strm0_tmp     ;
  reg [31:0] pe43_lane5_strm1 [0:4095];
  reg [31:0] pe43_lane5_strm1_tmp     ;
  reg [31:0] pe43_lane6_strm0 [0:4095];
  reg [31:0] pe43_lane6_strm0_tmp     ;
  reg [31:0] pe43_lane6_strm1 [0:4095];
  reg [31:0] pe43_lane6_strm1_tmp     ;
  reg [31:0] pe43_lane7_strm0 [0:4095];
  reg [31:0] pe43_lane7_strm0_tmp     ;
  reg [31:0] pe43_lane7_strm1 [0:4095];
  reg [31:0] pe43_lane7_strm1_tmp     ;
  reg [31:0] pe43_lane8_strm0 [0:4095];
  reg [31:0] pe43_lane8_strm0_tmp     ;
  reg [31:0] pe43_lane8_strm1 [0:4095];
  reg [31:0] pe43_lane8_strm1_tmp     ;
  reg [31:0] pe43_lane9_strm0 [0:4095];
  reg [31:0] pe43_lane9_strm0_tmp     ;
  reg [31:0] pe43_lane9_strm1 [0:4095];
  reg [31:0] pe43_lane9_strm1_tmp     ;
  reg [31:0] pe43_lane10_strm0 [0:4095];
  reg [31:0] pe43_lane10_strm0_tmp     ;
  reg [31:0] pe43_lane10_strm1 [0:4095];
  reg [31:0] pe43_lane10_strm1_tmp     ;
  reg [31:0] pe43_lane11_strm0 [0:4095];
  reg [31:0] pe43_lane11_strm0_tmp     ;
  reg [31:0] pe43_lane11_strm1 [0:4095];
  reg [31:0] pe43_lane11_strm1_tmp     ;
  reg [31:0] pe43_lane12_strm0 [0:4095];
  reg [31:0] pe43_lane12_strm0_tmp     ;
  reg [31:0] pe43_lane12_strm1 [0:4095];
  reg [31:0] pe43_lane12_strm1_tmp     ;
  reg [31:0] pe43_lane13_strm0 [0:4095];
  reg [31:0] pe43_lane13_strm0_tmp     ;
  reg [31:0] pe43_lane13_strm1 [0:4095];
  reg [31:0] pe43_lane13_strm1_tmp     ;
  reg [31:0] pe43_lane14_strm0 [0:4095];
  reg [31:0] pe43_lane14_strm0_tmp     ;
  reg [31:0] pe43_lane14_strm1 [0:4095];
  reg [31:0] pe43_lane14_strm1_tmp     ;
  reg [31:0] pe43_lane15_strm0 [0:4095];
  reg [31:0] pe43_lane15_strm0_tmp     ;
  reg [31:0] pe43_lane15_strm1 [0:4095];
  reg [31:0] pe43_lane15_strm1_tmp     ;
  reg [31:0] pe43_lane16_strm0 [0:4095];
  reg [31:0] pe43_lane16_strm0_tmp     ;
  reg [31:0] pe43_lane16_strm1 [0:4095];
  reg [31:0] pe43_lane16_strm1_tmp     ;
  reg [31:0] pe43_lane17_strm0 [0:4095];
  reg [31:0] pe43_lane17_strm0_tmp     ;
  reg [31:0] pe43_lane17_strm1 [0:4095];
  reg [31:0] pe43_lane17_strm1_tmp     ;
  reg [31:0] pe43_lane18_strm0 [0:4095];
  reg [31:0] pe43_lane18_strm0_tmp     ;
  reg [31:0] pe43_lane18_strm1 [0:4095];
  reg [31:0] pe43_lane18_strm1_tmp     ;
  reg [31:0] pe43_lane19_strm0 [0:4095];
  reg [31:0] pe43_lane19_strm0_tmp     ;
  reg [31:0] pe43_lane19_strm1 [0:4095];
  reg [31:0] pe43_lane19_strm1_tmp     ;
  reg [31:0] pe43_lane20_strm0 [0:4095];
  reg [31:0] pe43_lane20_strm0_tmp     ;
  reg [31:0] pe43_lane20_strm1 [0:4095];
  reg [31:0] pe43_lane20_strm1_tmp     ;
  reg [31:0] pe43_lane21_strm0 [0:4095];
  reg [31:0] pe43_lane21_strm0_tmp     ;
  reg [31:0] pe43_lane21_strm1 [0:4095];
  reg [31:0] pe43_lane21_strm1_tmp     ;
  reg [31:0] pe43_lane22_strm0 [0:4095];
  reg [31:0] pe43_lane22_strm0_tmp     ;
  reg [31:0] pe43_lane22_strm1 [0:4095];
  reg [31:0] pe43_lane22_strm1_tmp     ;
  reg [31:0] pe43_lane23_strm0 [0:4095];
  reg [31:0] pe43_lane23_strm0_tmp     ;
  reg [31:0] pe43_lane23_strm1 [0:4095];
  reg [31:0] pe43_lane23_strm1_tmp     ;
  reg [31:0] pe43_lane24_strm0 [0:4095];
  reg [31:0] pe43_lane24_strm0_tmp     ;
  reg [31:0] pe43_lane24_strm1 [0:4095];
  reg [31:0] pe43_lane24_strm1_tmp     ;
  reg [31:0] pe43_lane25_strm0 [0:4095];
  reg [31:0] pe43_lane25_strm0_tmp     ;
  reg [31:0] pe43_lane25_strm1 [0:4095];
  reg [31:0] pe43_lane25_strm1_tmp     ;
  reg [31:0] pe43_lane26_strm0 [0:4095];
  reg [31:0] pe43_lane26_strm0_tmp     ;
  reg [31:0] pe43_lane26_strm1 [0:4095];
  reg [31:0] pe43_lane26_strm1_tmp     ;
  reg [31:0] pe43_lane27_strm0 [0:4095];
  reg [31:0] pe43_lane27_strm0_tmp     ;
  reg [31:0] pe43_lane27_strm1 [0:4095];
  reg [31:0] pe43_lane27_strm1_tmp     ;
  reg [31:0] pe43_lane28_strm0 [0:4095];
  reg [31:0] pe43_lane28_strm0_tmp     ;
  reg [31:0] pe43_lane28_strm1 [0:4095];
  reg [31:0] pe43_lane28_strm1_tmp     ;
  reg [31:0] pe43_lane29_strm0 [0:4095];
  reg [31:0] pe43_lane29_strm0_tmp     ;
  reg [31:0] pe43_lane29_strm1 [0:4095];
  reg [31:0] pe43_lane29_strm1_tmp     ;
  reg [31:0] pe43_lane30_strm0 [0:4095];
  reg [31:0] pe43_lane30_strm0_tmp     ;
  reg [31:0] pe43_lane30_strm1 [0:4095];
  reg [31:0] pe43_lane30_strm1_tmp     ;
  reg [31:0] pe43_lane31_strm0 [0:4095];
  reg [31:0] pe43_lane31_strm0_tmp     ;
  reg [31:0] pe43_lane31_strm1 [0:4095];
  reg [31:0] pe43_lane31_strm1_tmp     ;
  reg [31:0] pe44_lane0_strm0 [0:4095];
  reg [31:0] pe44_lane0_strm0_tmp     ;
  reg [31:0] pe44_lane0_strm1 [0:4095];
  reg [31:0] pe44_lane0_strm1_tmp     ;
  reg [31:0] pe44_lane1_strm0 [0:4095];
  reg [31:0] pe44_lane1_strm0_tmp     ;
  reg [31:0] pe44_lane1_strm1 [0:4095];
  reg [31:0] pe44_lane1_strm1_tmp     ;
  reg [31:0] pe44_lane2_strm0 [0:4095];
  reg [31:0] pe44_lane2_strm0_tmp     ;
  reg [31:0] pe44_lane2_strm1 [0:4095];
  reg [31:0] pe44_lane2_strm1_tmp     ;
  reg [31:0] pe44_lane3_strm0 [0:4095];
  reg [31:0] pe44_lane3_strm0_tmp     ;
  reg [31:0] pe44_lane3_strm1 [0:4095];
  reg [31:0] pe44_lane3_strm1_tmp     ;
  reg [31:0] pe44_lane4_strm0 [0:4095];
  reg [31:0] pe44_lane4_strm0_tmp     ;
  reg [31:0] pe44_lane4_strm1 [0:4095];
  reg [31:0] pe44_lane4_strm1_tmp     ;
  reg [31:0] pe44_lane5_strm0 [0:4095];
  reg [31:0] pe44_lane5_strm0_tmp     ;
  reg [31:0] pe44_lane5_strm1 [0:4095];
  reg [31:0] pe44_lane5_strm1_tmp     ;
  reg [31:0] pe44_lane6_strm0 [0:4095];
  reg [31:0] pe44_lane6_strm0_tmp     ;
  reg [31:0] pe44_lane6_strm1 [0:4095];
  reg [31:0] pe44_lane6_strm1_tmp     ;
  reg [31:0] pe44_lane7_strm0 [0:4095];
  reg [31:0] pe44_lane7_strm0_tmp     ;
  reg [31:0] pe44_lane7_strm1 [0:4095];
  reg [31:0] pe44_lane7_strm1_tmp     ;
  reg [31:0] pe44_lane8_strm0 [0:4095];
  reg [31:0] pe44_lane8_strm0_tmp     ;
  reg [31:0] pe44_lane8_strm1 [0:4095];
  reg [31:0] pe44_lane8_strm1_tmp     ;
  reg [31:0] pe44_lane9_strm0 [0:4095];
  reg [31:0] pe44_lane9_strm0_tmp     ;
  reg [31:0] pe44_lane9_strm1 [0:4095];
  reg [31:0] pe44_lane9_strm1_tmp     ;
  reg [31:0] pe44_lane10_strm0 [0:4095];
  reg [31:0] pe44_lane10_strm0_tmp     ;
  reg [31:0] pe44_lane10_strm1 [0:4095];
  reg [31:0] pe44_lane10_strm1_tmp     ;
  reg [31:0] pe44_lane11_strm0 [0:4095];
  reg [31:0] pe44_lane11_strm0_tmp     ;
  reg [31:0] pe44_lane11_strm1 [0:4095];
  reg [31:0] pe44_lane11_strm1_tmp     ;
  reg [31:0] pe44_lane12_strm0 [0:4095];
  reg [31:0] pe44_lane12_strm0_tmp     ;
  reg [31:0] pe44_lane12_strm1 [0:4095];
  reg [31:0] pe44_lane12_strm1_tmp     ;
  reg [31:0] pe44_lane13_strm0 [0:4095];
  reg [31:0] pe44_lane13_strm0_tmp     ;
  reg [31:0] pe44_lane13_strm1 [0:4095];
  reg [31:0] pe44_lane13_strm1_tmp     ;
  reg [31:0] pe44_lane14_strm0 [0:4095];
  reg [31:0] pe44_lane14_strm0_tmp     ;
  reg [31:0] pe44_lane14_strm1 [0:4095];
  reg [31:0] pe44_lane14_strm1_tmp     ;
  reg [31:0] pe44_lane15_strm0 [0:4095];
  reg [31:0] pe44_lane15_strm0_tmp     ;
  reg [31:0] pe44_lane15_strm1 [0:4095];
  reg [31:0] pe44_lane15_strm1_tmp     ;
  reg [31:0] pe44_lane16_strm0 [0:4095];
  reg [31:0] pe44_lane16_strm0_tmp     ;
  reg [31:0] pe44_lane16_strm1 [0:4095];
  reg [31:0] pe44_lane16_strm1_tmp     ;
  reg [31:0] pe44_lane17_strm0 [0:4095];
  reg [31:0] pe44_lane17_strm0_tmp     ;
  reg [31:0] pe44_lane17_strm1 [0:4095];
  reg [31:0] pe44_lane17_strm1_tmp     ;
  reg [31:0] pe44_lane18_strm0 [0:4095];
  reg [31:0] pe44_lane18_strm0_tmp     ;
  reg [31:0] pe44_lane18_strm1 [0:4095];
  reg [31:0] pe44_lane18_strm1_tmp     ;
  reg [31:0] pe44_lane19_strm0 [0:4095];
  reg [31:0] pe44_lane19_strm0_tmp     ;
  reg [31:0] pe44_lane19_strm1 [0:4095];
  reg [31:0] pe44_lane19_strm1_tmp     ;
  reg [31:0] pe44_lane20_strm0 [0:4095];
  reg [31:0] pe44_lane20_strm0_tmp     ;
  reg [31:0] pe44_lane20_strm1 [0:4095];
  reg [31:0] pe44_lane20_strm1_tmp     ;
  reg [31:0] pe44_lane21_strm0 [0:4095];
  reg [31:0] pe44_lane21_strm0_tmp     ;
  reg [31:0] pe44_lane21_strm1 [0:4095];
  reg [31:0] pe44_lane21_strm1_tmp     ;
  reg [31:0] pe44_lane22_strm0 [0:4095];
  reg [31:0] pe44_lane22_strm0_tmp     ;
  reg [31:0] pe44_lane22_strm1 [0:4095];
  reg [31:0] pe44_lane22_strm1_tmp     ;
  reg [31:0] pe44_lane23_strm0 [0:4095];
  reg [31:0] pe44_lane23_strm0_tmp     ;
  reg [31:0] pe44_lane23_strm1 [0:4095];
  reg [31:0] pe44_lane23_strm1_tmp     ;
  reg [31:0] pe44_lane24_strm0 [0:4095];
  reg [31:0] pe44_lane24_strm0_tmp     ;
  reg [31:0] pe44_lane24_strm1 [0:4095];
  reg [31:0] pe44_lane24_strm1_tmp     ;
  reg [31:0] pe44_lane25_strm0 [0:4095];
  reg [31:0] pe44_lane25_strm0_tmp     ;
  reg [31:0] pe44_lane25_strm1 [0:4095];
  reg [31:0] pe44_lane25_strm1_tmp     ;
  reg [31:0] pe44_lane26_strm0 [0:4095];
  reg [31:0] pe44_lane26_strm0_tmp     ;
  reg [31:0] pe44_lane26_strm1 [0:4095];
  reg [31:0] pe44_lane26_strm1_tmp     ;
  reg [31:0] pe44_lane27_strm0 [0:4095];
  reg [31:0] pe44_lane27_strm0_tmp     ;
  reg [31:0] pe44_lane27_strm1 [0:4095];
  reg [31:0] pe44_lane27_strm1_tmp     ;
  reg [31:0] pe44_lane28_strm0 [0:4095];
  reg [31:0] pe44_lane28_strm0_tmp     ;
  reg [31:0] pe44_lane28_strm1 [0:4095];
  reg [31:0] pe44_lane28_strm1_tmp     ;
  reg [31:0] pe44_lane29_strm0 [0:4095];
  reg [31:0] pe44_lane29_strm0_tmp     ;
  reg [31:0] pe44_lane29_strm1 [0:4095];
  reg [31:0] pe44_lane29_strm1_tmp     ;
  reg [31:0] pe44_lane30_strm0 [0:4095];
  reg [31:0] pe44_lane30_strm0_tmp     ;
  reg [31:0] pe44_lane30_strm1 [0:4095];
  reg [31:0] pe44_lane30_strm1_tmp     ;
  reg [31:0] pe44_lane31_strm0 [0:4095];
  reg [31:0] pe44_lane31_strm0_tmp     ;
  reg [31:0] pe44_lane31_strm1 [0:4095];
  reg [31:0] pe44_lane31_strm1_tmp     ;
  reg [31:0] pe45_lane0_strm0 [0:4095];
  reg [31:0] pe45_lane0_strm0_tmp     ;
  reg [31:0] pe45_lane0_strm1 [0:4095];
  reg [31:0] pe45_lane0_strm1_tmp     ;
  reg [31:0] pe45_lane1_strm0 [0:4095];
  reg [31:0] pe45_lane1_strm0_tmp     ;
  reg [31:0] pe45_lane1_strm1 [0:4095];
  reg [31:0] pe45_lane1_strm1_tmp     ;
  reg [31:0] pe45_lane2_strm0 [0:4095];
  reg [31:0] pe45_lane2_strm0_tmp     ;
  reg [31:0] pe45_lane2_strm1 [0:4095];
  reg [31:0] pe45_lane2_strm1_tmp     ;
  reg [31:0] pe45_lane3_strm0 [0:4095];
  reg [31:0] pe45_lane3_strm0_tmp     ;
  reg [31:0] pe45_lane3_strm1 [0:4095];
  reg [31:0] pe45_lane3_strm1_tmp     ;
  reg [31:0] pe45_lane4_strm0 [0:4095];
  reg [31:0] pe45_lane4_strm0_tmp     ;
  reg [31:0] pe45_lane4_strm1 [0:4095];
  reg [31:0] pe45_lane4_strm1_tmp     ;
  reg [31:0] pe45_lane5_strm0 [0:4095];
  reg [31:0] pe45_lane5_strm0_tmp     ;
  reg [31:0] pe45_lane5_strm1 [0:4095];
  reg [31:0] pe45_lane5_strm1_tmp     ;
  reg [31:0] pe45_lane6_strm0 [0:4095];
  reg [31:0] pe45_lane6_strm0_tmp     ;
  reg [31:0] pe45_lane6_strm1 [0:4095];
  reg [31:0] pe45_lane6_strm1_tmp     ;
  reg [31:0] pe45_lane7_strm0 [0:4095];
  reg [31:0] pe45_lane7_strm0_tmp     ;
  reg [31:0] pe45_lane7_strm1 [0:4095];
  reg [31:0] pe45_lane7_strm1_tmp     ;
  reg [31:0] pe45_lane8_strm0 [0:4095];
  reg [31:0] pe45_lane8_strm0_tmp     ;
  reg [31:0] pe45_lane8_strm1 [0:4095];
  reg [31:0] pe45_lane8_strm1_tmp     ;
  reg [31:0] pe45_lane9_strm0 [0:4095];
  reg [31:0] pe45_lane9_strm0_tmp     ;
  reg [31:0] pe45_lane9_strm1 [0:4095];
  reg [31:0] pe45_lane9_strm1_tmp     ;
  reg [31:0] pe45_lane10_strm0 [0:4095];
  reg [31:0] pe45_lane10_strm0_tmp     ;
  reg [31:0] pe45_lane10_strm1 [0:4095];
  reg [31:0] pe45_lane10_strm1_tmp     ;
  reg [31:0] pe45_lane11_strm0 [0:4095];
  reg [31:0] pe45_lane11_strm0_tmp     ;
  reg [31:0] pe45_lane11_strm1 [0:4095];
  reg [31:0] pe45_lane11_strm1_tmp     ;
  reg [31:0] pe45_lane12_strm0 [0:4095];
  reg [31:0] pe45_lane12_strm0_tmp     ;
  reg [31:0] pe45_lane12_strm1 [0:4095];
  reg [31:0] pe45_lane12_strm1_tmp     ;
  reg [31:0] pe45_lane13_strm0 [0:4095];
  reg [31:0] pe45_lane13_strm0_tmp     ;
  reg [31:0] pe45_lane13_strm1 [0:4095];
  reg [31:0] pe45_lane13_strm1_tmp     ;
  reg [31:0] pe45_lane14_strm0 [0:4095];
  reg [31:0] pe45_lane14_strm0_tmp     ;
  reg [31:0] pe45_lane14_strm1 [0:4095];
  reg [31:0] pe45_lane14_strm1_tmp     ;
  reg [31:0] pe45_lane15_strm0 [0:4095];
  reg [31:0] pe45_lane15_strm0_tmp     ;
  reg [31:0] pe45_lane15_strm1 [0:4095];
  reg [31:0] pe45_lane15_strm1_tmp     ;
  reg [31:0] pe45_lane16_strm0 [0:4095];
  reg [31:0] pe45_lane16_strm0_tmp     ;
  reg [31:0] pe45_lane16_strm1 [0:4095];
  reg [31:0] pe45_lane16_strm1_tmp     ;
  reg [31:0] pe45_lane17_strm0 [0:4095];
  reg [31:0] pe45_lane17_strm0_tmp     ;
  reg [31:0] pe45_lane17_strm1 [0:4095];
  reg [31:0] pe45_lane17_strm1_tmp     ;
  reg [31:0] pe45_lane18_strm0 [0:4095];
  reg [31:0] pe45_lane18_strm0_tmp     ;
  reg [31:0] pe45_lane18_strm1 [0:4095];
  reg [31:0] pe45_lane18_strm1_tmp     ;
  reg [31:0] pe45_lane19_strm0 [0:4095];
  reg [31:0] pe45_lane19_strm0_tmp     ;
  reg [31:0] pe45_lane19_strm1 [0:4095];
  reg [31:0] pe45_lane19_strm1_tmp     ;
  reg [31:0] pe45_lane20_strm0 [0:4095];
  reg [31:0] pe45_lane20_strm0_tmp     ;
  reg [31:0] pe45_lane20_strm1 [0:4095];
  reg [31:0] pe45_lane20_strm1_tmp     ;
  reg [31:0] pe45_lane21_strm0 [0:4095];
  reg [31:0] pe45_lane21_strm0_tmp     ;
  reg [31:0] pe45_lane21_strm1 [0:4095];
  reg [31:0] pe45_lane21_strm1_tmp     ;
  reg [31:0] pe45_lane22_strm0 [0:4095];
  reg [31:0] pe45_lane22_strm0_tmp     ;
  reg [31:0] pe45_lane22_strm1 [0:4095];
  reg [31:0] pe45_lane22_strm1_tmp     ;
  reg [31:0] pe45_lane23_strm0 [0:4095];
  reg [31:0] pe45_lane23_strm0_tmp     ;
  reg [31:0] pe45_lane23_strm1 [0:4095];
  reg [31:0] pe45_lane23_strm1_tmp     ;
  reg [31:0] pe45_lane24_strm0 [0:4095];
  reg [31:0] pe45_lane24_strm0_tmp     ;
  reg [31:0] pe45_lane24_strm1 [0:4095];
  reg [31:0] pe45_lane24_strm1_tmp     ;
  reg [31:0] pe45_lane25_strm0 [0:4095];
  reg [31:0] pe45_lane25_strm0_tmp     ;
  reg [31:0] pe45_lane25_strm1 [0:4095];
  reg [31:0] pe45_lane25_strm1_tmp     ;
  reg [31:0] pe45_lane26_strm0 [0:4095];
  reg [31:0] pe45_lane26_strm0_tmp     ;
  reg [31:0] pe45_lane26_strm1 [0:4095];
  reg [31:0] pe45_lane26_strm1_tmp     ;
  reg [31:0] pe45_lane27_strm0 [0:4095];
  reg [31:0] pe45_lane27_strm0_tmp     ;
  reg [31:0] pe45_lane27_strm1 [0:4095];
  reg [31:0] pe45_lane27_strm1_tmp     ;
  reg [31:0] pe45_lane28_strm0 [0:4095];
  reg [31:0] pe45_lane28_strm0_tmp     ;
  reg [31:0] pe45_lane28_strm1 [0:4095];
  reg [31:0] pe45_lane28_strm1_tmp     ;
  reg [31:0] pe45_lane29_strm0 [0:4095];
  reg [31:0] pe45_lane29_strm0_tmp     ;
  reg [31:0] pe45_lane29_strm1 [0:4095];
  reg [31:0] pe45_lane29_strm1_tmp     ;
  reg [31:0] pe45_lane30_strm0 [0:4095];
  reg [31:0] pe45_lane30_strm0_tmp     ;
  reg [31:0] pe45_lane30_strm1 [0:4095];
  reg [31:0] pe45_lane30_strm1_tmp     ;
  reg [31:0] pe45_lane31_strm0 [0:4095];
  reg [31:0] pe45_lane31_strm0_tmp     ;
  reg [31:0] pe45_lane31_strm1 [0:4095];
  reg [31:0] pe45_lane31_strm1_tmp     ;
  reg [31:0] pe46_lane0_strm0 [0:4095];
  reg [31:0] pe46_lane0_strm0_tmp     ;
  reg [31:0] pe46_lane0_strm1 [0:4095];
  reg [31:0] pe46_lane0_strm1_tmp     ;
  reg [31:0] pe46_lane1_strm0 [0:4095];
  reg [31:0] pe46_lane1_strm0_tmp     ;
  reg [31:0] pe46_lane1_strm1 [0:4095];
  reg [31:0] pe46_lane1_strm1_tmp     ;
  reg [31:0] pe46_lane2_strm0 [0:4095];
  reg [31:0] pe46_lane2_strm0_tmp     ;
  reg [31:0] pe46_lane2_strm1 [0:4095];
  reg [31:0] pe46_lane2_strm1_tmp     ;
  reg [31:0] pe46_lane3_strm0 [0:4095];
  reg [31:0] pe46_lane3_strm0_tmp     ;
  reg [31:0] pe46_lane3_strm1 [0:4095];
  reg [31:0] pe46_lane3_strm1_tmp     ;
  reg [31:0] pe46_lane4_strm0 [0:4095];
  reg [31:0] pe46_lane4_strm0_tmp     ;
  reg [31:0] pe46_lane4_strm1 [0:4095];
  reg [31:0] pe46_lane4_strm1_tmp     ;
  reg [31:0] pe46_lane5_strm0 [0:4095];
  reg [31:0] pe46_lane5_strm0_tmp     ;
  reg [31:0] pe46_lane5_strm1 [0:4095];
  reg [31:0] pe46_lane5_strm1_tmp     ;
  reg [31:0] pe46_lane6_strm0 [0:4095];
  reg [31:0] pe46_lane6_strm0_tmp     ;
  reg [31:0] pe46_lane6_strm1 [0:4095];
  reg [31:0] pe46_lane6_strm1_tmp     ;
  reg [31:0] pe46_lane7_strm0 [0:4095];
  reg [31:0] pe46_lane7_strm0_tmp     ;
  reg [31:0] pe46_lane7_strm1 [0:4095];
  reg [31:0] pe46_lane7_strm1_tmp     ;
  reg [31:0] pe46_lane8_strm0 [0:4095];
  reg [31:0] pe46_lane8_strm0_tmp     ;
  reg [31:0] pe46_lane8_strm1 [0:4095];
  reg [31:0] pe46_lane8_strm1_tmp     ;
  reg [31:0] pe46_lane9_strm0 [0:4095];
  reg [31:0] pe46_lane9_strm0_tmp     ;
  reg [31:0] pe46_lane9_strm1 [0:4095];
  reg [31:0] pe46_lane9_strm1_tmp     ;
  reg [31:0] pe46_lane10_strm0 [0:4095];
  reg [31:0] pe46_lane10_strm0_tmp     ;
  reg [31:0] pe46_lane10_strm1 [0:4095];
  reg [31:0] pe46_lane10_strm1_tmp     ;
  reg [31:0] pe46_lane11_strm0 [0:4095];
  reg [31:0] pe46_lane11_strm0_tmp     ;
  reg [31:0] pe46_lane11_strm1 [0:4095];
  reg [31:0] pe46_lane11_strm1_tmp     ;
  reg [31:0] pe46_lane12_strm0 [0:4095];
  reg [31:0] pe46_lane12_strm0_tmp     ;
  reg [31:0] pe46_lane12_strm1 [0:4095];
  reg [31:0] pe46_lane12_strm1_tmp     ;
  reg [31:0] pe46_lane13_strm0 [0:4095];
  reg [31:0] pe46_lane13_strm0_tmp     ;
  reg [31:0] pe46_lane13_strm1 [0:4095];
  reg [31:0] pe46_lane13_strm1_tmp     ;
  reg [31:0] pe46_lane14_strm0 [0:4095];
  reg [31:0] pe46_lane14_strm0_tmp     ;
  reg [31:0] pe46_lane14_strm1 [0:4095];
  reg [31:0] pe46_lane14_strm1_tmp     ;
  reg [31:0] pe46_lane15_strm0 [0:4095];
  reg [31:0] pe46_lane15_strm0_tmp     ;
  reg [31:0] pe46_lane15_strm1 [0:4095];
  reg [31:0] pe46_lane15_strm1_tmp     ;
  reg [31:0] pe46_lane16_strm0 [0:4095];
  reg [31:0] pe46_lane16_strm0_tmp     ;
  reg [31:0] pe46_lane16_strm1 [0:4095];
  reg [31:0] pe46_lane16_strm1_tmp     ;
  reg [31:0] pe46_lane17_strm0 [0:4095];
  reg [31:0] pe46_lane17_strm0_tmp     ;
  reg [31:0] pe46_lane17_strm1 [0:4095];
  reg [31:0] pe46_lane17_strm1_tmp     ;
  reg [31:0] pe46_lane18_strm0 [0:4095];
  reg [31:0] pe46_lane18_strm0_tmp     ;
  reg [31:0] pe46_lane18_strm1 [0:4095];
  reg [31:0] pe46_lane18_strm1_tmp     ;
  reg [31:0] pe46_lane19_strm0 [0:4095];
  reg [31:0] pe46_lane19_strm0_tmp     ;
  reg [31:0] pe46_lane19_strm1 [0:4095];
  reg [31:0] pe46_lane19_strm1_tmp     ;
  reg [31:0] pe46_lane20_strm0 [0:4095];
  reg [31:0] pe46_lane20_strm0_tmp     ;
  reg [31:0] pe46_lane20_strm1 [0:4095];
  reg [31:0] pe46_lane20_strm1_tmp     ;
  reg [31:0] pe46_lane21_strm0 [0:4095];
  reg [31:0] pe46_lane21_strm0_tmp     ;
  reg [31:0] pe46_lane21_strm1 [0:4095];
  reg [31:0] pe46_lane21_strm1_tmp     ;
  reg [31:0] pe46_lane22_strm0 [0:4095];
  reg [31:0] pe46_lane22_strm0_tmp     ;
  reg [31:0] pe46_lane22_strm1 [0:4095];
  reg [31:0] pe46_lane22_strm1_tmp     ;
  reg [31:0] pe46_lane23_strm0 [0:4095];
  reg [31:0] pe46_lane23_strm0_tmp     ;
  reg [31:0] pe46_lane23_strm1 [0:4095];
  reg [31:0] pe46_lane23_strm1_tmp     ;
  reg [31:0] pe46_lane24_strm0 [0:4095];
  reg [31:0] pe46_lane24_strm0_tmp     ;
  reg [31:0] pe46_lane24_strm1 [0:4095];
  reg [31:0] pe46_lane24_strm1_tmp     ;
  reg [31:0] pe46_lane25_strm0 [0:4095];
  reg [31:0] pe46_lane25_strm0_tmp     ;
  reg [31:0] pe46_lane25_strm1 [0:4095];
  reg [31:0] pe46_lane25_strm1_tmp     ;
  reg [31:0] pe46_lane26_strm0 [0:4095];
  reg [31:0] pe46_lane26_strm0_tmp     ;
  reg [31:0] pe46_lane26_strm1 [0:4095];
  reg [31:0] pe46_lane26_strm1_tmp     ;
  reg [31:0] pe46_lane27_strm0 [0:4095];
  reg [31:0] pe46_lane27_strm0_tmp     ;
  reg [31:0] pe46_lane27_strm1 [0:4095];
  reg [31:0] pe46_lane27_strm1_tmp     ;
  reg [31:0] pe46_lane28_strm0 [0:4095];
  reg [31:0] pe46_lane28_strm0_tmp     ;
  reg [31:0] pe46_lane28_strm1 [0:4095];
  reg [31:0] pe46_lane28_strm1_tmp     ;
  reg [31:0] pe46_lane29_strm0 [0:4095];
  reg [31:0] pe46_lane29_strm0_tmp     ;
  reg [31:0] pe46_lane29_strm1 [0:4095];
  reg [31:0] pe46_lane29_strm1_tmp     ;
  reg [31:0] pe46_lane30_strm0 [0:4095];
  reg [31:0] pe46_lane30_strm0_tmp     ;
  reg [31:0] pe46_lane30_strm1 [0:4095];
  reg [31:0] pe46_lane30_strm1_tmp     ;
  reg [31:0] pe46_lane31_strm0 [0:4095];
  reg [31:0] pe46_lane31_strm0_tmp     ;
  reg [31:0] pe46_lane31_strm1 [0:4095];
  reg [31:0] pe46_lane31_strm1_tmp     ;
  reg [31:0] pe47_lane0_strm0 [0:4095];
  reg [31:0] pe47_lane0_strm0_tmp     ;
  reg [31:0] pe47_lane0_strm1 [0:4095];
  reg [31:0] pe47_lane0_strm1_tmp     ;
  reg [31:0] pe47_lane1_strm0 [0:4095];
  reg [31:0] pe47_lane1_strm0_tmp     ;
  reg [31:0] pe47_lane1_strm1 [0:4095];
  reg [31:0] pe47_lane1_strm1_tmp     ;
  reg [31:0] pe47_lane2_strm0 [0:4095];
  reg [31:0] pe47_lane2_strm0_tmp     ;
  reg [31:0] pe47_lane2_strm1 [0:4095];
  reg [31:0] pe47_lane2_strm1_tmp     ;
  reg [31:0] pe47_lane3_strm0 [0:4095];
  reg [31:0] pe47_lane3_strm0_tmp     ;
  reg [31:0] pe47_lane3_strm1 [0:4095];
  reg [31:0] pe47_lane3_strm1_tmp     ;
  reg [31:0] pe47_lane4_strm0 [0:4095];
  reg [31:0] pe47_lane4_strm0_tmp     ;
  reg [31:0] pe47_lane4_strm1 [0:4095];
  reg [31:0] pe47_lane4_strm1_tmp     ;
  reg [31:0] pe47_lane5_strm0 [0:4095];
  reg [31:0] pe47_lane5_strm0_tmp     ;
  reg [31:0] pe47_lane5_strm1 [0:4095];
  reg [31:0] pe47_lane5_strm1_tmp     ;
  reg [31:0] pe47_lane6_strm0 [0:4095];
  reg [31:0] pe47_lane6_strm0_tmp     ;
  reg [31:0] pe47_lane6_strm1 [0:4095];
  reg [31:0] pe47_lane6_strm1_tmp     ;
  reg [31:0] pe47_lane7_strm0 [0:4095];
  reg [31:0] pe47_lane7_strm0_tmp     ;
  reg [31:0] pe47_lane7_strm1 [0:4095];
  reg [31:0] pe47_lane7_strm1_tmp     ;
  reg [31:0] pe47_lane8_strm0 [0:4095];
  reg [31:0] pe47_lane8_strm0_tmp     ;
  reg [31:0] pe47_lane8_strm1 [0:4095];
  reg [31:0] pe47_lane8_strm1_tmp     ;
  reg [31:0] pe47_lane9_strm0 [0:4095];
  reg [31:0] pe47_lane9_strm0_tmp     ;
  reg [31:0] pe47_lane9_strm1 [0:4095];
  reg [31:0] pe47_lane9_strm1_tmp     ;
  reg [31:0] pe47_lane10_strm0 [0:4095];
  reg [31:0] pe47_lane10_strm0_tmp     ;
  reg [31:0] pe47_lane10_strm1 [0:4095];
  reg [31:0] pe47_lane10_strm1_tmp     ;
  reg [31:0] pe47_lane11_strm0 [0:4095];
  reg [31:0] pe47_lane11_strm0_tmp     ;
  reg [31:0] pe47_lane11_strm1 [0:4095];
  reg [31:0] pe47_lane11_strm1_tmp     ;
  reg [31:0] pe47_lane12_strm0 [0:4095];
  reg [31:0] pe47_lane12_strm0_tmp     ;
  reg [31:0] pe47_lane12_strm1 [0:4095];
  reg [31:0] pe47_lane12_strm1_tmp     ;
  reg [31:0] pe47_lane13_strm0 [0:4095];
  reg [31:0] pe47_lane13_strm0_tmp     ;
  reg [31:0] pe47_lane13_strm1 [0:4095];
  reg [31:0] pe47_lane13_strm1_tmp     ;
  reg [31:0] pe47_lane14_strm0 [0:4095];
  reg [31:0] pe47_lane14_strm0_tmp     ;
  reg [31:0] pe47_lane14_strm1 [0:4095];
  reg [31:0] pe47_lane14_strm1_tmp     ;
  reg [31:0] pe47_lane15_strm0 [0:4095];
  reg [31:0] pe47_lane15_strm0_tmp     ;
  reg [31:0] pe47_lane15_strm1 [0:4095];
  reg [31:0] pe47_lane15_strm1_tmp     ;
  reg [31:0] pe47_lane16_strm0 [0:4095];
  reg [31:0] pe47_lane16_strm0_tmp     ;
  reg [31:0] pe47_lane16_strm1 [0:4095];
  reg [31:0] pe47_lane16_strm1_tmp     ;
  reg [31:0] pe47_lane17_strm0 [0:4095];
  reg [31:0] pe47_lane17_strm0_tmp     ;
  reg [31:0] pe47_lane17_strm1 [0:4095];
  reg [31:0] pe47_lane17_strm1_tmp     ;
  reg [31:0] pe47_lane18_strm0 [0:4095];
  reg [31:0] pe47_lane18_strm0_tmp     ;
  reg [31:0] pe47_lane18_strm1 [0:4095];
  reg [31:0] pe47_lane18_strm1_tmp     ;
  reg [31:0] pe47_lane19_strm0 [0:4095];
  reg [31:0] pe47_lane19_strm0_tmp     ;
  reg [31:0] pe47_lane19_strm1 [0:4095];
  reg [31:0] pe47_lane19_strm1_tmp     ;
  reg [31:0] pe47_lane20_strm0 [0:4095];
  reg [31:0] pe47_lane20_strm0_tmp     ;
  reg [31:0] pe47_lane20_strm1 [0:4095];
  reg [31:0] pe47_lane20_strm1_tmp     ;
  reg [31:0] pe47_lane21_strm0 [0:4095];
  reg [31:0] pe47_lane21_strm0_tmp     ;
  reg [31:0] pe47_lane21_strm1 [0:4095];
  reg [31:0] pe47_lane21_strm1_tmp     ;
  reg [31:0] pe47_lane22_strm0 [0:4095];
  reg [31:0] pe47_lane22_strm0_tmp     ;
  reg [31:0] pe47_lane22_strm1 [0:4095];
  reg [31:0] pe47_lane22_strm1_tmp     ;
  reg [31:0] pe47_lane23_strm0 [0:4095];
  reg [31:0] pe47_lane23_strm0_tmp     ;
  reg [31:0] pe47_lane23_strm1 [0:4095];
  reg [31:0] pe47_lane23_strm1_tmp     ;
  reg [31:0] pe47_lane24_strm0 [0:4095];
  reg [31:0] pe47_lane24_strm0_tmp     ;
  reg [31:0] pe47_lane24_strm1 [0:4095];
  reg [31:0] pe47_lane24_strm1_tmp     ;
  reg [31:0] pe47_lane25_strm0 [0:4095];
  reg [31:0] pe47_lane25_strm0_tmp     ;
  reg [31:0] pe47_lane25_strm1 [0:4095];
  reg [31:0] pe47_lane25_strm1_tmp     ;
  reg [31:0] pe47_lane26_strm0 [0:4095];
  reg [31:0] pe47_lane26_strm0_tmp     ;
  reg [31:0] pe47_lane26_strm1 [0:4095];
  reg [31:0] pe47_lane26_strm1_tmp     ;
  reg [31:0] pe47_lane27_strm0 [0:4095];
  reg [31:0] pe47_lane27_strm0_tmp     ;
  reg [31:0] pe47_lane27_strm1 [0:4095];
  reg [31:0] pe47_lane27_strm1_tmp     ;
  reg [31:0] pe47_lane28_strm0 [0:4095];
  reg [31:0] pe47_lane28_strm0_tmp     ;
  reg [31:0] pe47_lane28_strm1 [0:4095];
  reg [31:0] pe47_lane28_strm1_tmp     ;
  reg [31:0] pe47_lane29_strm0 [0:4095];
  reg [31:0] pe47_lane29_strm0_tmp     ;
  reg [31:0] pe47_lane29_strm1 [0:4095];
  reg [31:0] pe47_lane29_strm1_tmp     ;
  reg [31:0] pe47_lane30_strm0 [0:4095];
  reg [31:0] pe47_lane30_strm0_tmp     ;
  reg [31:0] pe47_lane30_strm1 [0:4095];
  reg [31:0] pe47_lane30_strm1_tmp     ;
  reg [31:0] pe47_lane31_strm0 [0:4095];
  reg [31:0] pe47_lane31_strm0_tmp     ;
  reg [31:0] pe47_lane31_strm1 [0:4095];
  reg [31:0] pe47_lane31_strm1_tmp     ;
  reg [31:0] pe48_lane0_strm0 [0:4095];
  reg [31:0] pe48_lane0_strm0_tmp     ;
  reg [31:0] pe48_lane0_strm1 [0:4095];
  reg [31:0] pe48_lane0_strm1_tmp     ;
  reg [31:0] pe48_lane1_strm0 [0:4095];
  reg [31:0] pe48_lane1_strm0_tmp     ;
  reg [31:0] pe48_lane1_strm1 [0:4095];
  reg [31:0] pe48_lane1_strm1_tmp     ;
  reg [31:0] pe48_lane2_strm0 [0:4095];
  reg [31:0] pe48_lane2_strm0_tmp     ;
  reg [31:0] pe48_lane2_strm1 [0:4095];
  reg [31:0] pe48_lane2_strm1_tmp     ;
  reg [31:0] pe48_lane3_strm0 [0:4095];
  reg [31:0] pe48_lane3_strm0_tmp     ;
  reg [31:0] pe48_lane3_strm1 [0:4095];
  reg [31:0] pe48_lane3_strm1_tmp     ;
  reg [31:0] pe48_lane4_strm0 [0:4095];
  reg [31:0] pe48_lane4_strm0_tmp     ;
  reg [31:0] pe48_lane4_strm1 [0:4095];
  reg [31:0] pe48_lane4_strm1_tmp     ;
  reg [31:0] pe48_lane5_strm0 [0:4095];
  reg [31:0] pe48_lane5_strm0_tmp     ;
  reg [31:0] pe48_lane5_strm1 [0:4095];
  reg [31:0] pe48_lane5_strm1_tmp     ;
  reg [31:0] pe48_lane6_strm0 [0:4095];
  reg [31:0] pe48_lane6_strm0_tmp     ;
  reg [31:0] pe48_lane6_strm1 [0:4095];
  reg [31:0] pe48_lane6_strm1_tmp     ;
  reg [31:0] pe48_lane7_strm0 [0:4095];
  reg [31:0] pe48_lane7_strm0_tmp     ;
  reg [31:0] pe48_lane7_strm1 [0:4095];
  reg [31:0] pe48_lane7_strm1_tmp     ;
  reg [31:0] pe48_lane8_strm0 [0:4095];
  reg [31:0] pe48_lane8_strm0_tmp     ;
  reg [31:0] pe48_lane8_strm1 [0:4095];
  reg [31:0] pe48_lane8_strm1_tmp     ;
  reg [31:0] pe48_lane9_strm0 [0:4095];
  reg [31:0] pe48_lane9_strm0_tmp     ;
  reg [31:0] pe48_lane9_strm1 [0:4095];
  reg [31:0] pe48_lane9_strm1_tmp     ;
  reg [31:0] pe48_lane10_strm0 [0:4095];
  reg [31:0] pe48_lane10_strm0_tmp     ;
  reg [31:0] pe48_lane10_strm1 [0:4095];
  reg [31:0] pe48_lane10_strm1_tmp     ;
  reg [31:0] pe48_lane11_strm0 [0:4095];
  reg [31:0] pe48_lane11_strm0_tmp     ;
  reg [31:0] pe48_lane11_strm1 [0:4095];
  reg [31:0] pe48_lane11_strm1_tmp     ;
  reg [31:0] pe48_lane12_strm0 [0:4095];
  reg [31:0] pe48_lane12_strm0_tmp     ;
  reg [31:0] pe48_lane12_strm1 [0:4095];
  reg [31:0] pe48_lane12_strm1_tmp     ;
  reg [31:0] pe48_lane13_strm0 [0:4095];
  reg [31:0] pe48_lane13_strm0_tmp     ;
  reg [31:0] pe48_lane13_strm1 [0:4095];
  reg [31:0] pe48_lane13_strm1_tmp     ;
  reg [31:0] pe48_lane14_strm0 [0:4095];
  reg [31:0] pe48_lane14_strm0_tmp     ;
  reg [31:0] pe48_lane14_strm1 [0:4095];
  reg [31:0] pe48_lane14_strm1_tmp     ;
  reg [31:0] pe48_lane15_strm0 [0:4095];
  reg [31:0] pe48_lane15_strm0_tmp     ;
  reg [31:0] pe48_lane15_strm1 [0:4095];
  reg [31:0] pe48_lane15_strm1_tmp     ;
  reg [31:0] pe48_lane16_strm0 [0:4095];
  reg [31:0] pe48_lane16_strm0_tmp     ;
  reg [31:0] pe48_lane16_strm1 [0:4095];
  reg [31:0] pe48_lane16_strm1_tmp     ;
  reg [31:0] pe48_lane17_strm0 [0:4095];
  reg [31:0] pe48_lane17_strm0_tmp     ;
  reg [31:0] pe48_lane17_strm1 [0:4095];
  reg [31:0] pe48_lane17_strm1_tmp     ;
  reg [31:0] pe48_lane18_strm0 [0:4095];
  reg [31:0] pe48_lane18_strm0_tmp     ;
  reg [31:0] pe48_lane18_strm1 [0:4095];
  reg [31:0] pe48_lane18_strm1_tmp     ;
  reg [31:0] pe48_lane19_strm0 [0:4095];
  reg [31:0] pe48_lane19_strm0_tmp     ;
  reg [31:0] pe48_lane19_strm1 [0:4095];
  reg [31:0] pe48_lane19_strm1_tmp     ;
  reg [31:0] pe48_lane20_strm0 [0:4095];
  reg [31:0] pe48_lane20_strm0_tmp     ;
  reg [31:0] pe48_lane20_strm1 [0:4095];
  reg [31:0] pe48_lane20_strm1_tmp     ;
  reg [31:0] pe48_lane21_strm0 [0:4095];
  reg [31:0] pe48_lane21_strm0_tmp     ;
  reg [31:0] pe48_lane21_strm1 [0:4095];
  reg [31:0] pe48_lane21_strm1_tmp     ;
  reg [31:0] pe48_lane22_strm0 [0:4095];
  reg [31:0] pe48_lane22_strm0_tmp     ;
  reg [31:0] pe48_lane22_strm1 [0:4095];
  reg [31:0] pe48_lane22_strm1_tmp     ;
  reg [31:0] pe48_lane23_strm0 [0:4095];
  reg [31:0] pe48_lane23_strm0_tmp     ;
  reg [31:0] pe48_lane23_strm1 [0:4095];
  reg [31:0] pe48_lane23_strm1_tmp     ;
  reg [31:0] pe48_lane24_strm0 [0:4095];
  reg [31:0] pe48_lane24_strm0_tmp     ;
  reg [31:0] pe48_lane24_strm1 [0:4095];
  reg [31:0] pe48_lane24_strm1_tmp     ;
  reg [31:0] pe48_lane25_strm0 [0:4095];
  reg [31:0] pe48_lane25_strm0_tmp     ;
  reg [31:0] pe48_lane25_strm1 [0:4095];
  reg [31:0] pe48_lane25_strm1_tmp     ;
  reg [31:0] pe48_lane26_strm0 [0:4095];
  reg [31:0] pe48_lane26_strm0_tmp     ;
  reg [31:0] pe48_lane26_strm1 [0:4095];
  reg [31:0] pe48_lane26_strm1_tmp     ;
  reg [31:0] pe48_lane27_strm0 [0:4095];
  reg [31:0] pe48_lane27_strm0_tmp     ;
  reg [31:0] pe48_lane27_strm1 [0:4095];
  reg [31:0] pe48_lane27_strm1_tmp     ;
  reg [31:0] pe48_lane28_strm0 [0:4095];
  reg [31:0] pe48_lane28_strm0_tmp     ;
  reg [31:0] pe48_lane28_strm1 [0:4095];
  reg [31:0] pe48_lane28_strm1_tmp     ;
  reg [31:0] pe48_lane29_strm0 [0:4095];
  reg [31:0] pe48_lane29_strm0_tmp     ;
  reg [31:0] pe48_lane29_strm1 [0:4095];
  reg [31:0] pe48_lane29_strm1_tmp     ;
  reg [31:0] pe48_lane30_strm0 [0:4095];
  reg [31:0] pe48_lane30_strm0_tmp     ;
  reg [31:0] pe48_lane30_strm1 [0:4095];
  reg [31:0] pe48_lane30_strm1_tmp     ;
  reg [31:0] pe48_lane31_strm0 [0:4095];
  reg [31:0] pe48_lane31_strm0_tmp     ;
  reg [31:0] pe48_lane31_strm1 [0:4095];
  reg [31:0] pe48_lane31_strm1_tmp     ;
  reg [31:0] pe49_lane0_strm0 [0:4095];
  reg [31:0] pe49_lane0_strm0_tmp     ;
  reg [31:0] pe49_lane0_strm1 [0:4095];
  reg [31:0] pe49_lane0_strm1_tmp     ;
  reg [31:0] pe49_lane1_strm0 [0:4095];
  reg [31:0] pe49_lane1_strm0_tmp     ;
  reg [31:0] pe49_lane1_strm1 [0:4095];
  reg [31:0] pe49_lane1_strm1_tmp     ;
  reg [31:0] pe49_lane2_strm0 [0:4095];
  reg [31:0] pe49_lane2_strm0_tmp     ;
  reg [31:0] pe49_lane2_strm1 [0:4095];
  reg [31:0] pe49_lane2_strm1_tmp     ;
  reg [31:0] pe49_lane3_strm0 [0:4095];
  reg [31:0] pe49_lane3_strm0_tmp     ;
  reg [31:0] pe49_lane3_strm1 [0:4095];
  reg [31:0] pe49_lane3_strm1_tmp     ;
  reg [31:0] pe49_lane4_strm0 [0:4095];
  reg [31:0] pe49_lane4_strm0_tmp     ;
  reg [31:0] pe49_lane4_strm1 [0:4095];
  reg [31:0] pe49_lane4_strm1_tmp     ;
  reg [31:0] pe49_lane5_strm0 [0:4095];
  reg [31:0] pe49_lane5_strm0_tmp     ;
  reg [31:0] pe49_lane5_strm1 [0:4095];
  reg [31:0] pe49_lane5_strm1_tmp     ;
  reg [31:0] pe49_lane6_strm0 [0:4095];
  reg [31:0] pe49_lane6_strm0_tmp     ;
  reg [31:0] pe49_lane6_strm1 [0:4095];
  reg [31:0] pe49_lane6_strm1_tmp     ;
  reg [31:0] pe49_lane7_strm0 [0:4095];
  reg [31:0] pe49_lane7_strm0_tmp     ;
  reg [31:0] pe49_lane7_strm1 [0:4095];
  reg [31:0] pe49_lane7_strm1_tmp     ;
  reg [31:0] pe49_lane8_strm0 [0:4095];
  reg [31:0] pe49_lane8_strm0_tmp     ;
  reg [31:0] pe49_lane8_strm1 [0:4095];
  reg [31:0] pe49_lane8_strm1_tmp     ;
  reg [31:0] pe49_lane9_strm0 [0:4095];
  reg [31:0] pe49_lane9_strm0_tmp     ;
  reg [31:0] pe49_lane9_strm1 [0:4095];
  reg [31:0] pe49_lane9_strm1_tmp     ;
  reg [31:0] pe49_lane10_strm0 [0:4095];
  reg [31:0] pe49_lane10_strm0_tmp     ;
  reg [31:0] pe49_lane10_strm1 [0:4095];
  reg [31:0] pe49_lane10_strm1_tmp     ;
  reg [31:0] pe49_lane11_strm0 [0:4095];
  reg [31:0] pe49_lane11_strm0_tmp     ;
  reg [31:0] pe49_lane11_strm1 [0:4095];
  reg [31:0] pe49_lane11_strm1_tmp     ;
  reg [31:0] pe49_lane12_strm0 [0:4095];
  reg [31:0] pe49_lane12_strm0_tmp     ;
  reg [31:0] pe49_lane12_strm1 [0:4095];
  reg [31:0] pe49_lane12_strm1_tmp     ;
  reg [31:0] pe49_lane13_strm0 [0:4095];
  reg [31:0] pe49_lane13_strm0_tmp     ;
  reg [31:0] pe49_lane13_strm1 [0:4095];
  reg [31:0] pe49_lane13_strm1_tmp     ;
  reg [31:0] pe49_lane14_strm0 [0:4095];
  reg [31:0] pe49_lane14_strm0_tmp     ;
  reg [31:0] pe49_lane14_strm1 [0:4095];
  reg [31:0] pe49_lane14_strm1_tmp     ;
  reg [31:0] pe49_lane15_strm0 [0:4095];
  reg [31:0] pe49_lane15_strm0_tmp     ;
  reg [31:0] pe49_lane15_strm1 [0:4095];
  reg [31:0] pe49_lane15_strm1_tmp     ;
  reg [31:0] pe49_lane16_strm0 [0:4095];
  reg [31:0] pe49_lane16_strm0_tmp     ;
  reg [31:0] pe49_lane16_strm1 [0:4095];
  reg [31:0] pe49_lane16_strm1_tmp     ;
  reg [31:0] pe49_lane17_strm0 [0:4095];
  reg [31:0] pe49_lane17_strm0_tmp     ;
  reg [31:0] pe49_lane17_strm1 [0:4095];
  reg [31:0] pe49_lane17_strm1_tmp     ;
  reg [31:0] pe49_lane18_strm0 [0:4095];
  reg [31:0] pe49_lane18_strm0_tmp     ;
  reg [31:0] pe49_lane18_strm1 [0:4095];
  reg [31:0] pe49_lane18_strm1_tmp     ;
  reg [31:0] pe49_lane19_strm0 [0:4095];
  reg [31:0] pe49_lane19_strm0_tmp     ;
  reg [31:0] pe49_lane19_strm1 [0:4095];
  reg [31:0] pe49_lane19_strm1_tmp     ;
  reg [31:0] pe49_lane20_strm0 [0:4095];
  reg [31:0] pe49_lane20_strm0_tmp     ;
  reg [31:0] pe49_lane20_strm1 [0:4095];
  reg [31:0] pe49_lane20_strm1_tmp     ;
  reg [31:0] pe49_lane21_strm0 [0:4095];
  reg [31:0] pe49_lane21_strm0_tmp     ;
  reg [31:0] pe49_lane21_strm1 [0:4095];
  reg [31:0] pe49_lane21_strm1_tmp     ;
  reg [31:0] pe49_lane22_strm0 [0:4095];
  reg [31:0] pe49_lane22_strm0_tmp     ;
  reg [31:0] pe49_lane22_strm1 [0:4095];
  reg [31:0] pe49_lane22_strm1_tmp     ;
  reg [31:0] pe49_lane23_strm0 [0:4095];
  reg [31:0] pe49_lane23_strm0_tmp     ;
  reg [31:0] pe49_lane23_strm1 [0:4095];
  reg [31:0] pe49_lane23_strm1_tmp     ;
  reg [31:0] pe49_lane24_strm0 [0:4095];
  reg [31:0] pe49_lane24_strm0_tmp     ;
  reg [31:0] pe49_lane24_strm1 [0:4095];
  reg [31:0] pe49_lane24_strm1_tmp     ;
  reg [31:0] pe49_lane25_strm0 [0:4095];
  reg [31:0] pe49_lane25_strm0_tmp     ;
  reg [31:0] pe49_lane25_strm1 [0:4095];
  reg [31:0] pe49_lane25_strm1_tmp     ;
  reg [31:0] pe49_lane26_strm0 [0:4095];
  reg [31:0] pe49_lane26_strm0_tmp     ;
  reg [31:0] pe49_lane26_strm1 [0:4095];
  reg [31:0] pe49_lane26_strm1_tmp     ;
  reg [31:0] pe49_lane27_strm0 [0:4095];
  reg [31:0] pe49_lane27_strm0_tmp     ;
  reg [31:0] pe49_lane27_strm1 [0:4095];
  reg [31:0] pe49_lane27_strm1_tmp     ;
  reg [31:0] pe49_lane28_strm0 [0:4095];
  reg [31:0] pe49_lane28_strm0_tmp     ;
  reg [31:0] pe49_lane28_strm1 [0:4095];
  reg [31:0] pe49_lane28_strm1_tmp     ;
  reg [31:0] pe49_lane29_strm0 [0:4095];
  reg [31:0] pe49_lane29_strm0_tmp     ;
  reg [31:0] pe49_lane29_strm1 [0:4095];
  reg [31:0] pe49_lane29_strm1_tmp     ;
  reg [31:0] pe49_lane30_strm0 [0:4095];
  reg [31:0] pe49_lane30_strm0_tmp     ;
  reg [31:0] pe49_lane30_strm1 [0:4095];
  reg [31:0] pe49_lane30_strm1_tmp     ;
  reg [31:0] pe49_lane31_strm0 [0:4095];
  reg [31:0] pe49_lane31_strm0_tmp     ;
  reg [31:0] pe49_lane31_strm1 [0:4095];
  reg [31:0] pe49_lane31_strm1_tmp     ;
  reg [31:0] pe50_lane0_strm0 [0:4095];
  reg [31:0] pe50_lane0_strm0_tmp     ;
  reg [31:0] pe50_lane0_strm1 [0:4095];
  reg [31:0] pe50_lane0_strm1_tmp     ;
  reg [31:0] pe50_lane1_strm0 [0:4095];
  reg [31:0] pe50_lane1_strm0_tmp     ;
  reg [31:0] pe50_lane1_strm1 [0:4095];
  reg [31:0] pe50_lane1_strm1_tmp     ;
  reg [31:0] pe50_lane2_strm0 [0:4095];
  reg [31:0] pe50_lane2_strm0_tmp     ;
  reg [31:0] pe50_lane2_strm1 [0:4095];
  reg [31:0] pe50_lane2_strm1_tmp     ;
  reg [31:0] pe50_lane3_strm0 [0:4095];
  reg [31:0] pe50_lane3_strm0_tmp     ;
  reg [31:0] pe50_lane3_strm1 [0:4095];
  reg [31:0] pe50_lane3_strm1_tmp     ;
  reg [31:0] pe50_lane4_strm0 [0:4095];
  reg [31:0] pe50_lane4_strm0_tmp     ;
  reg [31:0] pe50_lane4_strm1 [0:4095];
  reg [31:0] pe50_lane4_strm1_tmp     ;
  reg [31:0] pe50_lane5_strm0 [0:4095];
  reg [31:0] pe50_lane5_strm0_tmp     ;
  reg [31:0] pe50_lane5_strm1 [0:4095];
  reg [31:0] pe50_lane5_strm1_tmp     ;
  reg [31:0] pe50_lane6_strm0 [0:4095];
  reg [31:0] pe50_lane6_strm0_tmp     ;
  reg [31:0] pe50_lane6_strm1 [0:4095];
  reg [31:0] pe50_lane6_strm1_tmp     ;
  reg [31:0] pe50_lane7_strm0 [0:4095];
  reg [31:0] pe50_lane7_strm0_tmp     ;
  reg [31:0] pe50_lane7_strm1 [0:4095];
  reg [31:0] pe50_lane7_strm1_tmp     ;
  reg [31:0] pe50_lane8_strm0 [0:4095];
  reg [31:0] pe50_lane8_strm0_tmp     ;
  reg [31:0] pe50_lane8_strm1 [0:4095];
  reg [31:0] pe50_lane8_strm1_tmp     ;
  reg [31:0] pe50_lane9_strm0 [0:4095];
  reg [31:0] pe50_lane9_strm0_tmp     ;
  reg [31:0] pe50_lane9_strm1 [0:4095];
  reg [31:0] pe50_lane9_strm1_tmp     ;
  reg [31:0] pe50_lane10_strm0 [0:4095];
  reg [31:0] pe50_lane10_strm0_tmp     ;
  reg [31:0] pe50_lane10_strm1 [0:4095];
  reg [31:0] pe50_lane10_strm1_tmp     ;
  reg [31:0] pe50_lane11_strm0 [0:4095];
  reg [31:0] pe50_lane11_strm0_tmp     ;
  reg [31:0] pe50_lane11_strm1 [0:4095];
  reg [31:0] pe50_lane11_strm1_tmp     ;
  reg [31:0] pe50_lane12_strm0 [0:4095];
  reg [31:0] pe50_lane12_strm0_tmp     ;
  reg [31:0] pe50_lane12_strm1 [0:4095];
  reg [31:0] pe50_lane12_strm1_tmp     ;
  reg [31:0] pe50_lane13_strm0 [0:4095];
  reg [31:0] pe50_lane13_strm0_tmp     ;
  reg [31:0] pe50_lane13_strm1 [0:4095];
  reg [31:0] pe50_lane13_strm1_tmp     ;
  reg [31:0] pe50_lane14_strm0 [0:4095];
  reg [31:0] pe50_lane14_strm0_tmp     ;
  reg [31:0] pe50_lane14_strm1 [0:4095];
  reg [31:0] pe50_lane14_strm1_tmp     ;
  reg [31:0] pe50_lane15_strm0 [0:4095];
  reg [31:0] pe50_lane15_strm0_tmp     ;
  reg [31:0] pe50_lane15_strm1 [0:4095];
  reg [31:0] pe50_lane15_strm1_tmp     ;
  reg [31:0] pe50_lane16_strm0 [0:4095];
  reg [31:0] pe50_lane16_strm0_tmp     ;
  reg [31:0] pe50_lane16_strm1 [0:4095];
  reg [31:0] pe50_lane16_strm1_tmp     ;
  reg [31:0] pe50_lane17_strm0 [0:4095];
  reg [31:0] pe50_lane17_strm0_tmp     ;
  reg [31:0] pe50_lane17_strm1 [0:4095];
  reg [31:0] pe50_lane17_strm1_tmp     ;
  reg [31:0] pe50_lane18_strm0 [0:4095];
  reg [31:0] pe50_lane18_strm0_tmp     ;
  reg [31:0] pe50_lane18_strm1 [0:4095];
  reg [31:0] pe50_lane18_strm1_tmp     ;
  reg [31:0] pe50_lane19_strm0 [0:4095];
  reg [31:0] pe50_lane19_strm0_tmp     ;
  reg [31:0] pe50_lane19_strm1 [0:4095];
  reg [31:0] pe50_lane19_strm1_tmp     ;
  reg [31:0] pe50_lane20_strm0 [0:4095];
  reg [31:0] pe50_lane20_strm0_tmp     ;
  reg [31:0] pe50_lane20_strm1 [0:4095];
  reg [31:0] pe50_lane20_strm1_tmp     ;
  reg [31:0] pe50_lane21_strm0 [0:4095];
  reg [31:0] pe50_lane21_strm0_tmp     ;
  reg [31:0] pe50_lane21_strm1 [0:4095];
  reg [31:0] pe50_lane21_strm1_tmp     ;
  reg [31:0] pe50_lane22_strm0 [0:4095];
  reg [31:0] pe50_lane22_strm0_tmp     ;
  reg [31:0] pe50_lane22_strm1 [0:4095];
  reg [31:0] pe50_lane22_strm1_tmp     ;
  reg [31:0] pe50_lane23_strm0 [0:4095];
  reg [31:0] pe50_lane23_strm0_tmp     ;
  reg [31:0] pe50_lane23_strm1 [0:4095];
  reg [31:0] pe50_lane23_strm1_tmp     ;
  reg [31:0] pe50_lane24_strm0 [0:4095];
  reg [31:0] pe50_lane24_strm0_tmp     ;
  reg [31:0] pe50_lane24_strm1 [0:4095];
  reg [31:0] pe50_lane24_strm1_tmp     ;
  reg [31:0] pe50_lane25_strm0 [0:4095];
  reg [31:0] pe50_lane25_strm0_tmp     ;
  reg [31:0] pe50_lane25_strm1 [0:4095];
  reg [31:0] pe50_lane25_strm1_tmp     ;
  reg [31:0] pe50_lane26_strm0 [0:4095];
  reg [31:0] pe50_lane26_strm0_tmp     ;
  reg [31:0] pe50_lane26_strm1 [0:4095];
  reg [31:0] pe50_lane26_strm1_tmp     ;
  reg [31:0] pe50_lane27_strm0 [0:4095];
  reg [31:0] pe50_lane27_strm0_tmp     ;
  reg [31:0] pe50_lane27_strm1 [0:4095];
  reg [31:0] pe50_lane27_strm1_tmp     ;
  reg [31:0] pe50_lane28_strm0 [0:4095];
  reg [31:0] pe50_lane28_strm0_tmp     ;
  reg [31:0] pe50_lane28_strm1 [0:4095];
  reg [31:0] pe50_lane28_strm1_tmp     ;
  reg [31:0] pe50_lane29_strm0 [0:4095];
  reg [31:0] pe50_lane29_strm0_tmp     ;
  reg [31:0] pe50_lane29_strm1 [0:4095];
  reg [31:0] pe50_lane29_strm1_tmp     ;
  reg [31:0] pe50_lane30_strm0 [0:4095];
  reg [31:0] pe50_lane30_strm0_tmp     ;
  reg [31:0] pe50_lane30_strm1 [0:4095];
  reg [31:0] pe50_lane30_strm1_tmp     ;
  reg [31:0] pe50_lane31_strm0 [0:4095];
  reg [31:0] pe50_lane31_strm0_tmp     ;
  reg [31:0] pe50_lane31_strm1 [0:4095];
  reg [31:0] pe50_lane31_strm1_tmp     ;
  reg [31:0] pe51_lane0_strm0 [0:4095];
  reg [31:0] pe51_lane0_strm0_tmp     ;
  reg [31:0] pe51_lane0_strm1 [0:4095];
  reg [31:0] pe51_lane0_strm1_tmp     ;
  reg [31:0] pe51_lane1_strm0 [0:4095];
  reg [31:0] pe51_lane1_strm0_tmp     ;
  reg [31:0] pe51_lane1_strm1 [0:4095];
  reg [31:0] pe51_lane1_strm1_tmp     ;
  reg [31:0] pe51_lane2_strm0 [0:4095];
  reg [31:0] pe51_lane2_strm0_tmp     ;
  reg [31:0] pe51_lane2_strm1 [0:4095];
  reg [31:0] pe51_lane2_strm1_tmp     ;
  reg [31:0] pe51_lane3_strm0 [0:4095];
  reg [31:0] pe51_lane3_strm0_tmp     ;
  reg [31:0] pe51_lane3_strm1 [0:4095];
  reg [31:0] pe51_lane3_strm1_tmp     ;
  reg [31:0] pe51_lane4_strm0 [0:4095];
  reg [31:0] pe51_lane4_strm0_tmp     ;
  reg [31:0] pe51_lane4_strm1 [0:4095];
  reg [31:0] pe51_lane4_strm1_tmp     ;
  reg [31:0] pe51_lane5_strm0 [0:4095];
  reg [31:0] pe51_lane5_strm0_tmp     ;
  reg [31:0] pe51_lane5_strm1 [0:4095];
  reg [31:0] pe51_lane5_strm1_tmp     ;
  reg [31:0] pe51_lane6_strm0 [0:4095];
  reg [31:0] pe51_lane6_strm0_tmp     ;
  reg [31:0] pe51_lane6_strm1 [0:4095];
  reg [31:0] pe51_lane6_strm1_tmp     ;
  reg [31:0] pe51_lane7_strm0 [0:4095];
  reg [31:0] pe51_lane7_strm0_tmp     ;
  reg [31:0] pe51_lane7_strm1 [0:4095];
  reg [31:0] pe51_lane7_strm1_tmp     ;
  reg [31:0] pe51_lane8_strm0 [0:4095];
  reg [31:0] pe51_lane8_strm0_tmp     ;
  reg [31:0] pe51_lane8_strm1 [0:4095];
  reg [31:0] pe51_lane8_strm1_tmp     ;
  reg [31:0] pe51_lane9_strm0 [0:4095];
  reg [31:0] pe51_lane9_strm0_tmp     ;
  reg [31:0] pe51_lane9_strm1 [0:4095];
  reg [31:0] pe51_lane9_strm1_tmp     ;
  reg [31:0] pe51_lane10_strm0 [0:4095];
  reg [31:0] pe51_lane10_strm0_tmp     ;
  reg [31:0] pe51_lane10_strm1 [0:4095];
  reg [31:0] pe51_lane10_strm1_tmp     ;
  reg [31:0] pe51_lane11_strm0 [0:4095];
  reg [31:0] pe51_lane11_strm0_tmp     ;
  reg [31:0] pe51_lane11_strm1 [0:4095];
  reg [31:0] pe51_lane11_strm1_tmp     ;
  reg [31:0] pe51_lane12_strm0 [0:4095];
  reg [31:0] pe51_lane12_strm0_tmp     ;
  reg [31:0] pe51_lane12_strm1 [0:4095];
  reg [31:0] pe51_lane12_strm1_tmp     ;
  reg [31:0] pe51_lane13_strm0 [0:4095];
  reg [31:0] pe51_lane13_strm0_tmp     ;
  reg [31:0] pe51_lane13_strm1 [0:4095];
  reg [31:0] pe51_lane13_strm1_tmp     ;
  reg [31:0] pe51_lane14_strm0 [0:4095];
  reg [31:0] pe51_lane14_strm0_tmp     ;
  reg [31:0] pe51_lane14_strm1 [0:4095];
  reg [31:0] pe51_lane14_strm1_tmp     ;
  reg [31:0] pe51_lane15_strm0 [0:4095];
  reg [31:0] pe51_lane15_strm0_tmp     ;
  reg [31:0] pe51_lane15_strm1 [0:4095];
  reg [31:0] pe51_lane15_strm1_tmp     ;
  reg [31:0] pe51_lane16_strm0 [0:4095];
  reg [31:0] pe51_lane16_strm0_tmp     ;
  reg [31:0] pe51_lane16_strm1 [0:4095];
  reg [31:0] pe51_lane16_strm1_tmp     ;
  reg [31:0] pe51_lane17_strm0 [0:4095];
  reg [31:0] pe51_lane17_strm0_tmp     ;
  reg [31:0] pe51_lane17_strm1 [0:4095];
  reg [31:0] pe51_lane17_strm1_tmp     ;
  reg [31:0] pe51_lane18_strm0 [0:4095];
  reg [31:0] pe51_lane18_strm0_tmp     ;
  reg [31:0] pe51_lane18_strm1 [0:4095];
  reg [31:0] pe51_lane18_strm1_tmp     ;
  reg [31:0] pe51_lane19_strm0 [0:4095];
  reg [31:0] pe51_lane19_strm0_tmp     ;
  reg [31:0] pe51_lane19_strm1 [0:4095];
  reg [31:0] pe51_lane19_strm1_tmp     ;
  reg [31:0] pe51_lane20_strm0 [0:4095];
  reg [31:0] pe51_lane20_strm0_tmp     ;
  reg [31:0] pe51_lane20_strm1 [0:4095];
  reg [31:0] pe51_lane20_strm1_tmp     ;
  reg [31:0] pe51_lane21_strm0 [0:4095];
  reg [31:0] pe51_lane21_strm0_tmp     ;
  reg [31:0] pe51_lane21_strm1 [0:4095];
  reg [31:0] pe51_lane21_strm1_tmp     ;
  reg [31:0] pe51_lane22_strm0 [0:4095];
  reg [31:0] pe51_lane22_strm0_tmp     ;
  reg [31:0] pe51_lane22_strm1 [0:4095];
  reg [31:0] pe51_lane22_strm1_tmp     ;
  reg [31:0] pe51_lane23_strm0 [0:4095];
  reg [31:0] pe51_lane23_strm0_tmp     ;
  reg [31:0] pe51_lane23_strm1 [0:4095];
  reg [31:0] pe51_lane23_strm1_tmp     ;
  reg [31:0] pe51_lane24_strm0 [0:4095];
  reg [31:0] pe51_lane24_strm0_tmp     ;
  reg [31:0] pe51_lane24_strm1 [0:4095];
  reg [31:0] pe51_lane24_strm1_tmp     ;
  reg [31:0] pe51_lane25_strm0 [0:4095];
  reg [31:0] pe51_lane25_strm0_tmp     ;
  reg [31:0] pe51_lane25_strm1 [0:4095];
  reg [31:0] pe51_lane25_strm1_tmp     ;
  reg [31:0] pe51_lane26_strm0 [0:4095];
  reg [31:0] pe51_lane26_strm0_tmp     ;
  reg [31:0] pe51_lane26_strm1 [0:4095];
  reg [31:0] pe51_lane26_strm1_tmp     ;
  reg [31:0] pe51_lane27_strm0 [0:4095];
  reg [31:0] pe51_lane27_strm0_tmp     ;
  reg [31:0] pe51_lane27_strm1 [0:4095];
  reg [31:0] pe51_lane27_strm1_tmp     ;
  reg [31:0] pe51_lane28_strm0 [0:4095];
  reg [31:0] pe51_lane28_strm0_tmp     ;
  reg [31:0] pe51_lane28_strm1 [0:4095];
  reg [31:0] pe51_lane28_strm1_tmp     ;
  reg [31:0] pe51_lane29_strm0 [0:4095];
  reg [31:0] pe51_lane29_strm0_tmp     ;
  reg [31:0] pe51_lane29_strm1 [0:4095];
  reg [31:0] pe51_lane29_strm1_tmp     ;
  reg [31:0] pe51_lane30_strm0 [0:4095];
  reg [31:0] pe51_lane30_strm0_tmp     ;
  reg [31:0] pe51_lane30_strm1 [0:4095];
  reg [31:0] pe51_lane30_strm1_tmp     ;
  reg [31:0] pe51_lane31_strm0 [0:4095];
  reg [31:0] pe51_lane31_strm0_tmp     ;
  reg [31:0] pe51_lane31_strm1 [0:4095];
  reg [31:0] pe51_lane31_strm1_tmp     ;
  reg [31:0] pe52_lane0_strm0 [0:4095];
  reg [31:0] pe52_lane0_strm0_tmp     ;
  reg [31:0] pe52_lane0_strm1 [0:4095];
  reg [31:0] pe52_lane0_strm1_tmp     ;
  reg [31:0] pe52_lane1_strm0 [0:4095];
  reg [31:0] pe52_lane1_strm0_tmp     ;
  reg [31:0] pe52_lane1_strm1 [0:4095];
  reg [31:0] pe52_lane1_strm1_tmp     ;
  reg [31:0] pe52_lane2_strm0 [0:4095];
  reg [31:0] pe52_lane2_strm0_tmp     ;
  reg [31:0] pe52_lane2_strm1 [0:4095];
  reg [31:0] pe52_lane2_strm1_tmp     ;
  reg [31:0] pe52_lane3_strm0 [0:4095];
  reg [31:0] pe52_lane3_strm0_tmp     ;
  reg [31:0] pe52_lane3_strm1 [0:4095];
  reg [31:0] pe52_lane3_strm1_tmp     ;
  reg [31:0] pe52_lane4_strm0 [0:4095];
  reg [31:0] pe52_lane4_strm0_tmp     ;
  reg [31:0] pe52_lane4_strm1 [0:4095];
  reg [31:0] pe52_lane4_strm1_tmp     ;
  reg [31:0] pe52_lane5_strm0 [0:4095];
  reg [31:0] pe52_lane5_strm0_tmp     ;
  reg [31:0] pe52_lane5_strm1 [0:4095];
  reg [31:0] pe52_lane5_strm1_tmp     ;
  reg [31:0] pe52_lane6_strm0 [0:4095];
  reg [31:0] pe52_lane6_strm0_tmp     ;
  reg [31:0] pe52_lane6_strm1 [0:4095];
  reg [31:0] pe52_lane6_strm1_tmp     ;
  reg [31:0] pe52_lane7_strm0 [0:4095];
  reg [31:0] pe52_lane7_strm0_tmp     ;
  reg [31:0] pe52_lane7_strm1 [0:4095];
  reg [31:0] pe52_lane7_strm1_tmp     ;
  reg [31:0] pe52_lane8_strm0 [0:4095];
  reg [31:0] pe52_lane8_strm0_tmp     ;
  reg [31:0] pe52_lane8_strm1 [0:4095];
  reg [31:0] pe52_lane8_strm1_tmp     ;
  reg [31:0] pe52_lane9_strm0 [0:4095];
  reg [31:0] pe52_lane9_strm0_tmp     ;
  reg [31:0] pe52_lane9_strm1 [0:4095];
  reg [31:0] pe52_lane9_strm1_tmp     ;
  reg [31:0] pe52_lane10_strm0 [0:4095];
  reg [31:0] pe52_lane10_strm0_tmp     ;
  reg [31:0] pe52_lane10_strm1 [0:4095];
  reg [31:0] pe52_lane10_strm1_tmp     ;
  reg [31:0] pe52_lane11_strm0 [0:4095];
  reg [31:0] pe52_lane11_strm0_tmp     ;
  reg [31:0] pe52_lane11_strm1 [0:4095];
  reg [31:0] pe52_lane11_strm1_tmp     ;
  reg [31:0] pe52_lane12_strm0 [0:4095];
  reg [31:0] pe52_lane12_strm0_tmp     ;
  reg [31:0] pe52_lane12_strm1 [0:4095];
  reg [31:0] pe52_lane12_strm1_tmp     ;
  reg [31:0] pe52_lane13_strm0 [0:4095];
  reg [31:0] pe52_lane13_strm0_tmp     ;
  reg [31:0] pe52_lane13_strm1 [0:4095];
  reg [31:0] pe52_lane13_strm1_tmp     ;
  reg [31:0] pe52_lane14_strm0 [0:4095];
  reg [31:0] pe52_lane14_strm0_tmp     ;
  reg [31:0] pe52_lane14_strm1 [0:4095];
  reg [31:0] pe52_lane14_strm1_tmp     ;
  reg [31:0] pe52_lane15_strm0 [0:4095];
  reg [31:0] pe52_lane15_strm0_tmp     ;
  reg [31:0] pe52_lane15_strm1 [0:4095];
  reg [31:0] pe52_lane15_strm1_tmp     ;
  reg [31:0] pe52_lane16_strm0 [0:4095];
  reg [31:0] pe52_lane16_strm0_tmp     ;
  reg [31:0] pe52_lane16_strm1 [0:4095];
  reg [31:0] pe52_lane16_strm1_tmp     ;
  reg [31:0] pe52_lane17_strm0 [0:4095];
  reg [31:0] pe52_lane17_strm0_tmp     ;
  reg [31:0] pe52_lane17_strm1 [0:4095];
  reg [31:0] pe52_lane17_strm1_tmp     ;
  reg [31:0] pe52_lane18_strm0 [0:4095];
  reg [31:0] pe52_lane18_strm0_tmp     ;
  reg [31:0] pe52_lane18_strm1 [0:4095];
  reg [31:0] pe52_lane18_strm1_tmp     ;
  reg [31:0] pe52_lane19_strm0 [0:4095];
  reg [31:0] pe52_lane19_strm0_tmp     ;
  reg [31:0] pe52_lane19_strm1 [0:4095];
  reg [31:0] pe52_lane19_strm1_tmp     ;
  reg [31:0] pe52_lane20_strm0 [0:4095];
  reg [31:0] pe52_lane20_strm0_tmp     ;
  reg [31:0] pe52_lane20_strm1 [0:4095];
  reg [31:0] pe52_lane20_strm1_tmp     ;
  reg [31:0] pe52_lane21_strm0 [0:4095];
  reg [31:0] pe52_lane21_strm0_tmp     ;
  reg [31:0] pe52_lane21_strm1 [0:4095];
  reg [31:0] pe52_lane21_strm1_tmp     ;
  reg [31:0] pe52_lane22_strm0 [0:4095];
  reg [31:0] pe52_lane22_strm0_tmp     ;
  reg [31:0] pe52_lane22_strm1 [0:4095];
  reg [31:0] pe52_lane22_strm1_tmp     ;
  reg [31:0] pe52_lane23_strm0 [0:4095];
  reg [31:0] pe52_lane23_strm0_tmp     ;
  reg [31:0] pe52_lane23_strm1 [0:4095];
  reg [31:0] pe52_lane23_strm1_tmp     ;
  reg [31:0] pe52_lane24_strm0 [0:4095];
  reg [31:0] pe52_lane24_strm0_tmp     ;
  reg [31:0] pe52_lane24_strm1 [0:4095];
  reg [31:0] pe52_lane24_strm1_tmp     ;
  reg [31:0] pe52_lane25_strm0 [0:4095];
  reg [31:0] pe52_lane25_strm0_tmp     ;
  reg [31:0] pe52_lane25_strm1 [0:4095];
  reg [31:0] pe52_lane25_strm1_tmp     ;
  reg [31:0] pe52_lane26_strm0 [0:4095];
  reg [31:0] pe52_lane26_strm0_tmp     ;
  reg [31:0] pe52_lane26_strm1 [0:4095];
  reg [31:0] pe52_lane26_strm1_tmp     ;
  reg [31:0] pe52_lane27_strm0 [0:4095];
  reg [31:0] pe52_lane27_strm0_tmp     ;
  reg [31:0] pe52_lane27_strm1 [0:4095];
  reg [31:0] pe52_lane27_strm1_tmp     ;
  reg [31:0] pe52_lane28_strm0 [0:4095];
  reg [31:0] pe52_lane28_strm0_tmp     ;
  reg [31:0] pe52_lane28_strm1 [0:4095];
  reg [31:0] pe52_lane28_strm1_tmp     ;
  reg [31:0] pe52_lane29_strm0 [0:4095];
  reg [31:0] pe52_lane29_strm0_tmp     ;
  reg [31:0] pe52_lane29_strm1 [0:4095];
  reg [31:0] pe52_lane29_strm1_tmp     ;
  reg [31:0] pe52_lane30_strm0 [0:4095];
  reg [31:0] pe52_lane30_strm0_tmp     ;
  reg [31:0] pe52_lane30_strm1 [0:4095];
  reg [31:0] pe52_lane30_strm1_tmp     ;
  reg [31:0] pe52_lane31_strm0 [0:4095];
  reg [31:0] pe52_lane31_strm0_tmp     ;
  reg [31:0] pe52_lane31_strm1 [0:4095];
  reg [31:0] pe52_lane31_strm1_tmp     ;
  reg [31:0] pe53_lane0_strm0 [0:4095];
  reg [31:0] pe53_lane0_strm0_tmp     ;
  reg [31:0] pe53_lane0_strm1 [0:4095];
  reg [31:0] pe53_lane0_strm1_tmp     ;
  reg [31:0] pe53_lane1_strm0 [0:4095];
  reg [31:0] pe53_lane1_strm0_tmp     ;
  reg [31:0] pe53_lane1_strm1 [0:4095];
  reg [31:0] pe53_lane1_strm1_tmp     ;
  reg [31:0] pe53_lane2_strm0 [0:4095];
  reg [31:0] pe53_lane2_strm0_tmp     ;
  reg [31:0] pe53_lane2_strm1 [0:4095];
  reg [31:0] pe53_lane2_strm1_tmp     ;
  reg [31:0] pe53_lane3_strm0 [0:4095];
  reg [31:0] pe53_lane3_strm0_tmp     ;
  reg [31:0] pe53_lane3_strm1 [0:4095];
  reg [31:0] pe53_lane3_strm1_tmp     ;
  reg [31:0] pe53_lane4_strm0 [0:4095];
  reg [31:0] pe53_lane4_strm0_tmp     ;
  reg [31:0] pe53_lane4_strm1 [0:4095];
  reg [31:0] pe53_lane4_strm1_tmp     ;
  reg [31:0] pe53_lane5_strm0 [0:4095];
  reg [31:0] pe53_lane5_strm0_tmp     ;
  reg [31:0] pe53_lane5_strm1 [0:4095];
  reg [31:0] pe53_lane5_strm1_tmp     ;
  reg [31:0] pe53_lane6_strm0 [0:4095];
  reg [31:0] pe53_lane6_strm0_tmp     ;
  reg [31:0] pe53_lane6_strm1 [0:4095];
  reg [31:0] pe53_lane6_strm1_tmp     ;
  reg [31:0] pe53_lane7_strm0 [0:4095];
  reg [31:0] pe53_lane7_strm0_tmp     ;
  reg [31:0] pe53_lane7_strm1 [0:4095];
  reg [31:0] pe53_lane7_strm1_tmp     ;
  reg [31:0] pe53_lane8_strm0 [0:4095];
  reg [31:0] pe53_lane8_strm0_tmp     ;
  reg [31:0] pe53_lane8_strm1 [0:4095];
  reg [31:0] pe53_lane8_strm1_tmp     ;
  reg [31:0] pe53_lane9_strm0 [0:4095];
  reg [31:0] pe53_lane9_strm0_tmp     ;
  reg [31:0] pe53_lane9_strm1 [0:4095];
  reg [31:0] pe53_lane9_strm1_tmp     ;
  reg [31:0] pe53_lane10_strm0 [0:4095];
  reg [31:0] pe53_lane10_strm0_tmp     ;
  reg [31:0] pe53_lane10_strm1 [0:4095];
  reg [31:0] pe53_lane10_strm1_tmp     ;
  reg [31:0] pe53_lane11_strm0 [0:4095];
  reg [31:0] pe53_lane11_strm0_tmp     ;
  reg [31:0] pe53_lane11_strm1 [0:4095];
  reg [31:0] pe53_lane11_strm1_tmp     ;
  reg [31:0] pe53_lane12_strm0 [0:4095];
  reg [31:0] pe53_lane12_strm0_tmp     ;
  reg [31:0] pe53_lane12_strm1 [0:4095];
  reg [31:0] pe53_lane12_strm1_tmp     ;
  reg [31:0] pe53_lane13_strm0 [0:4095];
  reg [31:0] pe53_lane13_strm0_tmp     ;
  reg [31:0] pe53_lane13_strm1 [0:4095];
  reg [31:0] pe53_lane13_strm1_tmp     ;
  reg [31:0] pe53_lane14_strm0 [0:4095];
  reg [31:0] pe53_lane14_strm0_tmp     ;
  reg [31:0] pe53_lane14_strm1 [0:4095];
  reg [31:0] pe53_lane14_strm1_tmp     ;
  reg [31:0] pe53_lane15_strm0 [0:4095];
  reg [31:0] pe53_lane15_strm0_tmp     ;
  reg [31:0] pe53_lane15_strm1 [0:4095];
  reg [31:0] pe53_lane15_strm1_tmp     ;
  reg [31:0] pe53_lane16_strm0 [0:4095];
  reg [31:0] pe53_lane16_strm0_tmp     ;
  reg [31:0] pe53_lane16_strm1 [0:4095];
  reg [31:0] pe53_lane16_strm1_tmp     ;
  reg [31:0] pe53_lane17_strm0 [0:4095];
  reg [31:0] pe53_lane17_strm0_tmp     ;
  reg [31:0] pe53_lane17_strm1 [0:4095];
  reg [31:0] pe53_lane17_strm1_tmp     ;
  reg [31:0] pe53_lane18_strm0 [0:4095];
  reg [31:0] pe53_lane18_strm0_tmp     ;
  reg [31:0] pe53_lane18_strm1 [0:4095];
  reg [31:0] pe53_lane18_strm1_tmp     ;
  reg [31:0] pe53_lane19_strm0 [0:4095];
  reg [31:0] pe53_lane19_strm0_tmp     ;
  reg [31:0] pe53_lane19_strm1 [0:4095];
  reg [31:0] pe53_lane19_strm1_tmp     ;
  reg [31:0] pe53_lane20_strm0 [0:4095];
  reg [31:0] pe53_lane20_strm0_tmp     ;
  reg [31:0] pe53_lane20_strm1 [0:4095];
  reg [31:0] pe53_lane20_strm1_tmp     ;
  reg [31:0] pe53_lane21_strm0 [0:4095];
  reg [31:0] pe53_lane21_strm0_tmp     ;
  reg [31:0] pe53_lane21_strm1 [0:4095];
  reg [31:0] pe53_lane21_strm1_tmp     ;
  reg [31:0] pe53_lane22_strm0 [0:4095];
  reg [31:0] pe53_lane22_strm0_tmp     ;
  reg [31:0] pe53_lane22_strm1 [0:4095];
  reg [31:0] pe53_lane22_strm1_tmp     ;
  reg [31:0] pe53_lane23_strm0 [0:4095];
  reg [31:0] pe53_lane23_strm0_tmp     ;
  reg [31:0] pe53_lane23_strm1 [0:4095];
  reg [31:0] pe53_lane23_strm1_tmp     ;
  reg [31:0] pe53_lane24_strm0 [0:4095];
  reg [31:0] pe53_lane24_strm0_tmp     ;
  reg [31:0] pe53_lane24_strm1 [0:4095];
  reg [31:0] pe53_lane24_strm1_tmp     ;
  reg [31:0] pe53_lane25_strm0 [0:4095];
  reg [31:0] pe53_lane25_strm0_tmp     ;
  reg [31:0] pe53_lane25_strm1 [0:4095];
  reg [31:0] pe53_lane25_strm1_tmp     ;
  reg [31:0] pe53_lane26_strm0 [0:4095];
  reg [31:0] pe53_lane26_strm0_tmp     ;
  reg [31:0] pe53_lane26_strm1 [0:4095];
  reg [31:0] pe53_lane26_strm1_tmp     ;
  reg [31:0] pe53_lane27_strm0 [0:4095];
  reg [31:0] pe53_lane27_strm0_tmp     ;
  reg [31:0] pe53_lane27_strm1 [0:4095];
  reg [31:0] pe53_lane27_strm1_tmp     ;
  reg [31:0] pe53_lane28_strm0 [0:4095];
  reg [31:0] pe53_lane28_strm0_tmp     ;
  reg [31:0] pe53_lane28_strm1 [0:4095];
  reg [31:0] pe53_lane28_strm1_tmp     ;
  reg [31:0] pe53_lane29_strm0 [0:4095];
  reg [31:0] pe53_lane29_strm0_tmp     ;
  reg [31:0] pe53_lane29_strm1 [0:4095];
  reg [31:0] pe53_lane29_strm1_tmp     ;
  reg [31:0] pe53_lane30_strm0 [0:4095];
  reg [31:0] pe53_lane30_strm0_tmp     ;
  reg [31:0] pe53_lane30_strm1 [0:4095];
  reg [31:0] pe53_lane30_strm1_tmp     ;
  reg [31:0] pe53_lane31_strm0 [0:4095];
  reg [31:0] pe53_lane31_strm0_tmp     ;
  reg [31:0] pe53_lane31_strm1 [0:4095];
  reg [31:0] pe53_lane31_strm1_tmp     ;
  reg [31:0] pe54_lane0_strm0 [0:4095];
  reg [31:0] pe54_lane0_strm0_tmp     ;
  reg [31:0] pe54_lane0_strm1 [0:4095];
  reg [31:0] pe54_lane0_strm1_tmp     ;
  reg [31:0] pe54_lane1_strm0 [0:4095];
  reg [31:0] pe54_lane1_strm0_tmp     ;
  reg [31:0] pe54_lane1_strm1 [0:4095];
  reg [31:0] pe54_lane1_strm1_tmp     ;
  reg [31:0] pe54_lane2_strm0 [0:4095];
  reg [31:0] pe54_lane2_strm0_tmp     ;
  reg [31:0] pe54_lane2_strm1 [0:4095];
  reg [31:0] pe54_lane2_strm1_tmp     ;
  reg [31:0] pe54_lane3_strm0 [0:4095];
  reg [31:0] pe54_lane3_strm0_tmp     ;
  reg [31:0] pe54_lane3_strm1 [0:4095];
  reg [31:0] pe54_lane3_strm1_tmp     ;
  reg [31:0] pe54_lane4_strm0 [0:4095];
  reg [31:0] pe54_lane4_strm0_tmp     ;
  reg [31:0] pe54_lane4_strm1 [0:4095];
  reg [31:0] pe54_lane4_strm1_tmp     ;
  reg [31:0] pe54_lane5_strm0 [0:4095];
  reg [31:0] pe54_lane5_strm0_tmp     ;
  reg [31:0] pe54_lane5_strm1 [0:4095];
  reg [31:0] pe54_lane5_strm1_tmp     ;
  reg [31:0] pe54_lane6_strm0 [0:4095];
  reg [31:0] pe54_lane6_strm0_tmp     ;
  reg [31:0] pe54_lane6_strm1 [0:4095];
  reg [31:0] pe54_lane6_strm1_tmp     ;
  reg [31:0] pe54_lane7_strm0 [0:4095];
  reg [31:0] pe54_lane7_strm0_tmp     ;
  reg [31:0] pe54_lane7_strm1 [0:4095];
  reg [31:0] pe54_lane7_strm1_tmp     ;
  reg [31:0] pe54_lane8_strm0 [0:4095];
  reg [31:0] pe54_lane8_strm0_tmp     ;
  reg [31:0] pe54_lane8_strm1 [0:4095];
  reg [31:0] pe54_lane8_strm1_tmp     ;
  reg [31:0] pe54_lane9_strm0 [0:4095];
  reg [31:0] pe54_lane9_strm0_tmp     ;
  reg [31:0] pe54_lane9_strm1 [0:4095];
  reg [31:0] pe54_lane9_strm1_tmp     ;
  reg [31:0] pe54_lane10_strm0 [0:4095];
  reg [31:0] pe54_lane10_strm0_tmp     ;
  reg [31:0] pe54_lane10_strm1 [0:4095];
  reg [31:0] pe54_lane10_strm1_tmp     ;
  reg [31:0] pe54_lane11_strm0 [0:4095];
  reg [31:0] pe54_lane11_strm0_tmp     ;
  reg [31:0] pe54_lane11_strm1 [0:4095];
  reg [31:0] pe54_lane11_strm1_tmp     ;
  reg [31:0] pe54_lane12_strm0 [0:4095];
  reg [31:0] pe54_lane12_strm0_tmp     ;
  reg [31:0] pe54_lane12_strm1 [0:4095];
  reg [31:0] pe54_lane12_strm1_tmp     ;
  reg [31:0] pe54_lane13_strm0 [0:4095];
  reg [31:0] pe54_lane13_strm0_tmp     ;
  reg [31:0] pe54_lane13_strm1 [0:4095];
  reg [31:0] pe54_lane13_strm1_tmp     ;
  reg [31:0] pe54_lane14_strm0 [0:4095];
  reg [31:0] pe54_lane14_strm0_tmp     ;
  reg [31:0] pe54_lane14_strm1 [0:4095];
  reg [31:0] pe54_lane14_strm1_tmp     ;
  reg [31:0] pe54_lane15_strm0 [0:4095];
  reg [31:0] pe54_lane15_strm0_tmp     ;
  reg [31:0] pe54_lane15_strm1 [0:4095];
  reg [31:0] pe54_lane15_strm1_tmp     ;
  reg [31:0] pe54_lane16_strm0 [0:4095];
  reg [31:0] pe54_lane16_strm0_tmp     ;
  reg [31:0] pe54_lane16_strm1 [0:4095];
  reg [31:0] pe54_lane16_strm1_tmp     ;
  reg [31:0] pe54_lane17_strm0 [0:4095];
  reg [31:0] pe54_lane17_strm0_tmp     ;
  reg [31:0] pe54_lane17_strm1 [0:4095];
  reg [31:0] pe54_lane17_strm1_tmp     ;
  reg [31:0] pe54_lane18_strm0 [0:4095];
  reg [31:0] pe54_lane18_strm0_tmp     ;
  reg [31:0] pe54_lane18_strm1 [0:4095];
  reg [31:0] pe54_lane18_strm1_tmp     ;
  reg [31:0] pe54_lane19_strm0 [0:4095];
  reg [31:0] pe54_lane19_strm0_tmp     ;
  reg [31:0] pe54_lane19_strm1 [0:4095];
  reg [31:0] pe54_lane19_strm1_tmp     ;
  reg [31:0] pe54_lane20_strm0 [0:4095];
  reg [31:0] pe54_lane20_strm0_tmp     ;
  reg [31:0] pe54_lane20_strm1 [0:4095];
  reg [31:0] pe54_lane20_strm1_tmp     ;
  reg [31:0] pe54_lane21_strm0 [0:4095];
  reg [31:0] pe54_lane21_strm0_tmp     ;
  reg [31:0] pe54_lane21_strm1 [0:4095];
  reg [31:0] pe54_lane21_strm1_tmp     ;
  reg [31:0] pe54_lane22_strm0 [0:4095];
  reg [31:0] pe54_lane22_strm0_tmp     ;
  reg [31:0] pe54_lane22_strm1 [0:4095];
  reg [31:0] pe54_lane22_strm1_tmp     ;
  reg [31:0] pe54_lane23_strm0 [0:4095];
  reg [31:0] pe54_lane23_strm0_tmp     ;
  reg [31:0] pe54_lane23_strm1 [0:4095];
  reg [31:0] pe54_lane23_strm1_tmp     ;
  reg [31:0] pe54_lane24_strm0 [0:4095];
  reg [31:0] pe54_lane24_strm0_tmp     ;
  reg [31:0] pe54_lane24_strm1 [0:4095];
  reg [31:0] pe54_lane24_strm1_tmp     ;
  reg [31:0] pe54_lane25_strm0 [0:4095];
  reg [31:0] pe54_lane25_strm0_tmp     ;
  reg [31:0] pe54_lane25_strm1 [0:4095];
  reg [31:0] pe54_lane25_strm1_tmp     ;
  reg [31:0] pe54_lane26_strm0 [0:4095];
  reg [31:0] pe54_lane26_strm0_tmp     ;
  reg [31:0] pe54_lane26_strm1 [0:4095];
  reg [31:0] pe54_lane26_strm1_tmp     ;
  reg [31:0] pe54_lane27_strm0 [0:4095];
  reg [31:0] pe54_lane27_strm0_tmp     ;
  reg [31:0] pe54_lane27_strm1 [0:4095];
  reg [31:0] pe54_lane27_strm1_tmp     ;
  reg [31:0] pe54_lane28_strm0 [0:4095];
  reg [31:0] pe54_lane28_strm0_tmp     ;
  reg [31:0] pe54_lane28_strm1 [0:4095];
  reg [31:0] pe54_lane28_strm1_tmp     ;
  reg [31:0] pe54_lane29_strm0 [0:4095];
  reg [31:0] pe54_lane29_strm0_tmp     ;
  reg [31:0] pe54_lane29_strm1 [0:4095];
  reg [31:0] pe54_lane29_strm1_tmp     ;
  reg [31:0] pe54_lane30_strm0 [0:4095];
  reg [31:0] pe54_lane30_strm0_tmp     ;
  reg [31:0] pe54_lane30_strm1 [0:4095];
  reg [31:0] pe54_lane30_strm1_tmp     ;
  reg [31:0] pe54_lane31_strm0 [0:4095];
  reg [31:0] pe54_lane31_strm0_tmp     ;
  reg [31:0] pe54_lane31_strm1 [0:4095];
  reg [31:0] pe54_lane31_strm1_tmp     ;
  reg [31:0] pe55_lane0_strm0 [0:4095];
  reg [31:0] pe55_lane0_strm0_tmp     ;
  reg [31:0] pe55_lane0_strm1 [0:4095];
  reg [31:0] pe55_lane0_strm1_tmp     ;
  reg [31:0] pe55_lane1_strm0 [0:4095];
  reg [31:0] pe55_lane1_strm0_tmp     ;
  reg [31:0] pe55_lane1_strm1 [0:4095];
  reg [31:0] pe55_lane1_strm1_tmp     ;
  reg [31:0] pe55_lane2_strm0 [0:4095];
  reg [31:0] pe55_lane2_strm0_tmp     ;
  reg [31:0] pe55_lane2_strm1 [0:4095];
  reg [31:0] pe55_lane2_strm1_tmp     ;
  reg [31:0] pe55_lane3_strm0 [0:4095];
  reg [31:0] pe55_lane3_strm0_tmp     ;
  reg [31:0] pe55_lane3_strm1 [0:4095];
  reg [31:0] pe55_lane3_strm1_tmp     ;
  reg [31:0] pe55_lane4_strm0 [0:4095];
  reg [31:0] pe55_lane4_strm0_tmp     ;
  reg [31:0] pe55_lane4_strm1 [0:4095];
  reg [31:0] pe55_lane4_strm1_tmp     ;
  reg [31:0] pe55_lane5_strm0 [0:4095];
  reg [31:0] pe55_lane5_strm0_tmp     ;
  reg [31:0] pe55_lane5_strm1 [0:4095];
  reg [31:0] pe55_lane5_strm1_tmp     ;
  reg [31:0] pe55_lane6_strm0 [0:4095];
  reg [31:0] pe55_lane6_strm0_tmp     ;
  reg [31:0] pe55_lane6_strm1 [0:4095];
  reg [31:0] pe55_lane6_strm1_tmp     ;
  reg [31:0] pe55_lane7_strm0 [0:4095];
  reg [31:0] pe55_lane7_strm0_tmp     ;
  reg [31:0] pe55_lane7_strm1 [0:4095];
  reg [31:0] pe55_lane7_strm1_tmp     ;
  reg [31:0] pe55_lane8_strm0 [0:4095];
  reg [31:0] pe55_lane8_strm0_tmp     ;
  reg [31:0] pe55_lane8_strm1 [0:4095];
  reg [31:0] pe55_lane8_strm1_tmp     ;
  reg [31:0] pe55_lane9_strm0 [0:4095];
  reg [31:0] pe55_lane9_strm0_tmp     ;
  reg [31:0] pe55_lane9_strm1 [0:4095];
  reg [31:0] pe55_lane9_strm1_tmp     ;
  reg [31:0] pe55_lane10_strm0 [0:4095];
  reg [31:0] pe55_lane10_strm0_tmp     ;
  reg [31:0] pe55_lane10_strm1 [0:4095];
  reg [31:0] pe55_lane10_strm1_tmp     ;
  reg [31:0] pe55_lane11_strm0 [0:4095];
  reg [31:0] pe55_lane11_strm0_tmp     ;
  reg [31:0] pe55_lane11_strm1 [0:4095];
  reg [31:0] pe55_lane11_strm1_tmp     ;
  reg [31:0] pe55_lane12_strm0 [0:4095];
  reg [31:0] pe55_lane12_strm0_tmp     ;
  reg [31:0] pe55_lane12_strm1 [0:4095];
  reg [31:0] pe55_lane12_strm1_tmp     ;
  reg [31:0] pe55_lane13_strm0 [0:4095];
  reg [31:0] pe55_lane13_strm0_tmp     ;
  reg [31:0] pe55_lane13_strm1 [0:4095];
  reg [31:0] pe55_lane13_strm1_tmp     ;
  reg [31:0] pe55_lane14_strm0 [0:4095];
  reg [31:0] pe55_lane14_strm0_tmp     ;
  reg [31:0] pe55_lane14_strm1 [0:4095];
  reg [31:0] pe55_lane14_strm1_tmp     ;
  reg [31:0] pe55_lane15_strm0 [0:4095];
  reg [31:0] pe55_lane15_strm0_tmp     ;
  reg [31:0] pe55_lane15_strm1 [0:4095];
  reg [31:0] pe55_lane15_strm1_tmp     ;
  reg [31:0] pe55_lane16_strm0 [0:4095];
  reg [31:0] pe55_lane16_strm0_tmp     ;
  reg [31:0] pe55_lane16_strm1 [0:4095];
  reg [31:0] pe55_lane16_strm1_tmp     ;
  reg [31:0] pe55_lane17_strm0 [0:4095];
  reg [31:0] pe55_lane17_strm0_tmp     ;
  reg [31:0] pe55_lane17_strm1 [0:4095];
  reg [31:0] pe55_lane17_strm1_tmp     ;
  reg [31:0] pe55_lane18_strm0 [0:4095];
  reg [31:0] pe55_lane18_strm0_tmp     ;
  reg [31:0] pe55_lane18_strm1 [0:4095];
  reg [31:0] pe55_lane18_strm1_tmp     ;
  reg [31:0] pe55_lane19_strm0 [0:4095];
  reg [31:0] pe55_lane19_strm0_tmp     ;
  reg [31:0] pe55_lane19_strm1 [0:4095];
  reg [31:0] pe55_lane19_strm1_tmp     ;
  reg [31:0] pe55_lane20_strm0 [0:4095];
  reg [31:0] pe55_lane20_strm0_tmp     ;
  reg [31:0] pe55_lane20_strm1 [0:4095];
  reg [31:0] pe55_lane20_strm1_tmp     ;
  reg [31:0] pe55_lane21_strm0 [0:4095];
  reg [31:0] pe55_lane21_strm0_tmp     ;
  reg [31:0] pe55_lane21_strm1 [0:4095];
  reg [31:0] pe55_lane21_strm1_tmp     ;
  reg [31:0] pe55_lane22_strm0 [0:4095];
  reg [31:0] pe55_lane22_strm0_tmp     ;
  reg [31:0] pe55_lane22_strm1 [0:4095];
  reg [31:0] pe55_lane22_strm1_tmp     ;
  reg [31:0] pe55_lane23_strm0 [0:4095];
  reg [31:0] pe55_lane23_strm0_tmp     ;
  reg [31:0] pe55_lane23_strm1 [0:4095];
  reg [31:0] pe55_lane23_strm1_tmp     ;
  reg [31:0] pe55_lane24_strm0 [0:4095];
  reg [31:0] pe55_lane24_strm0_tmp     ;
  reg [31:0] pe55_lane24_strm1 [0:4095];
  reg [31:0] pe55_lane24_strm1_tmp     ;
  reg [31:0] pe55_lane25_strm0 [0:4095];
  reg [31:0] pe55_lane25_strm0_tmp     ;
  reg [31:0] pe55_lane25_strm1 [0:4095];
  reg [31:0] pe55_lane25_strm1_tmp     ;
  reg [31:0] pe55_lane26_strm0 [0:4095];
  reg [31:0] pe55_lane26_strm0_tmp     ;
  reg [31:0] pe55_lane26_strm1 [0:4095];
  reg [31:0] pe55_lane26_strm1_tmp     ;
  reg [31:0] pe55_lane27_strm0 [0:4095];
  reg [31:0] pe55_lane27_strm0_tmp     ;
  reg [31:0] pe55_lane27_strm1 [0:4095];
  reg [31:0] pe55_lane27_strm1_tmp     ;
  reg [31:0] pe55_lane28_strm0 [0:4095];
  reg [31:0] pe55_lane28_strm0_tmp     ;
  reg [31:0] pe55_lane28_strm1 [0:4095];
  reg [31:0] pe55_lane28_strm1_tmp     ;
  reg [31:0] pe55_lane29_strm0 [0:4095];
  reg [31:0] pe55_lane29_strm0_tmp     ;
  reg [31:0] pe55_lane29_strm1 [0:4095];
  reg [31:0] pe55_lane29_strm1_tmp     ;
  reg [31:0] pe55_lane30_strm0 [0:4095];
  reg [31:0] pe55_lane30_strm0_tmp     ;
  reg [31:0] pe55_lane30_strm1 [0:4095];
  reg [31:0] pe55_lane30_strm1_tmp     ;
  reg [31:0] pe55_lane31_strm0 [0:4095];
  reg [31:0] pe55_lane31_strm0_tmp     ;
  reg [31:0] pe55_lane31_strm1 [0:4095];
  reg [31:0] pe55_lane31_strm1_tmp     ;
  reg [31:0] pe56_lane0_strm0 [0:4095];
  reg [31:0] pe56_lane0_strm0_tmp     ;
  reg [31:0] pe56_lane0_strm1 [0:4095];
  reg [31:0] pe56_lane0_strm1_tmp     ;
  reg [31:0] pe56_lane1_strm0 [0:4095];
  reg [31:0] pe56_lane1_strm0_tmp     ;
  reg [31:0] pe56_lane1_strm1 [0:4095];
  reg [31:0] pe56_lane1_strm1_tmp     ;
  reg [31:0] pe56_lane2_strm0 [0:4095];
  reg [31:0] pe56_lane2_strm0_tmp     ;
  reg [31:0] pe56_lane2_strm1 [0:4095];
  reg [31:0] pe56_lane2_strm1_tmp     ;
  reg [31:0] pe56_lane3_strm0 [0:4095];
  reg [31:0] pe56_lane3_strm0_tmp     ;
  reg [31:0] pe56_lane3_strm1 [0:4095];
  reg [31:0] pe56_lane3_strm1_tmp     ;
  reg [31:0] pe56_lane4_strm0 [0:4095];
  reg [31:0] pe56_lane4_strm0_tmp     ;
  reg [31:0] pe56_lane4_strm1 [0:4095];
  reg [31:0] pe56_lane4_strm1_tmp     ;
  reg [31:0] pe56_lane5_strm0 [0:4095];
  reg [31:0] pe56_lane5_strm0_tmp     ;
  reg [31:0] pe56_lane5_strm1 [0:4095];
  reg [31:0] pe56_lane5_strm1_tmp     ;
  reg [31:0] pe56_lane6_strm0 [0:4095];
  reg [31:0] pe56_lane6_strm0_tmp     ;
  reg [31:0] pe56_lane6_strm1 [0:4095];
  reg [31:0] pe56_lane6_strm1_tmp     ;
  reg [31:0] pe56_lane7_strm0 [0:4095];
  reg [31:0] pe56_lane7_strm0_tmp     ;
  reg [31:0] pe56_lane7_strm1 [0:4095];
  reg [31:0] pe56_lane7_strm1_tmp     ;
  reg [31:0] pe56_lane8_strm0 [0:4095];
  reg [31:0] pe56_lane8_strm0_tmp     ;
  reg [31:0] pe56_lane8_strm1 [0:4095];
  reg [31:0] pe56_lane8_strm1_tmp     ;
  reg [31:0] pe56_lane9_strm0 [0:4095];
  reg [31:0] pe56_lane9_strm0_tmp     ;
  reg [31:0] pe56_lane9_strm1 [0:4095];
  reg [31:0] pe56_lane9_strm1_tmp     ;
  reg [31:0] pe56_lane10_strm0 [0:4095];
  reg [31:0] pe56_lane10_strm0_tmp     ;
  reg [31:0] pe56_lane10_strm1 [0:4095];
  reg [31:0] pe56_lane10_strm1_tmp     ;
  reg [31:0] pe56_lane11_strm0 [0:4095];
  reg [31:0] pe56_lane11_strm0_tmp     ;
  reg [31:0] pe56_lane11_strm1 [0:4095];
  reg [31:0] pe56_lane11_strm1_tmp     ;
  reg [31:0] pe56_lane12_strm0 [0:4095];
  reg [31:0] pe56_lane12_strm0_tmp     ;
  reg [31:0] pe56_lane12_strm1 [0:4095];
  reg [31:0] pe56_lane12_strm1_tmp     ;
  reg [31:0] pe56_lane13_strm0 [0:4095];
  reg [31:0] pe56_lane13_strm0_tmp     ;
  reg [31:0] pe56_lane13_strm1 [0:4095];
  reg [31:0] pe56_lane13_strm1_tmp     ;
  reg [31:0] pe56_lane14_strm0 [0:4095];
  reg [31:0] pe56_lane14_strm0_tmp     ;
  reg [31:0] pe56_lane14_strm1 [0:4095];
  reg [31:0] pe56_lane14_strm1_tmp     ;
  reg [31:0] pe56_lane15_strm0 [0:4095];
  reg [31:0] pe56_lane15_strm0_tmp     ;
  reg [31:0] pe56_lane15_strm1 [0:4095];
  reg [31:0] pe56_lane15_strm1_tmp     ;
  reg [31:0] pe56_lane16_strm0 [0:4095];
  reg [31:0] pe56_lane16_strm0_tmp     ;
  reg [31:0] pe56_lane16_strm1 [0:4095];
  reg [31:0] pe56_lane16_strm1_tmp     ;
  reg [31:0] pe56_lane17_strm0 [0:4095];
  reg [31:0] pe56_lane17_strm0_tmp     ;
  reg [31:0] pe56_lane17_strm1 [0:4095];
  reg [31:0] pe56_lane17_strm1_tmp     ;
  reg [31:0] pe56_lane18_strm0 [0:4095];
  reg [31:0] pe56_lane18_strm0_tmp     ;
  reg [31:0] pe56_lane18_strm1 [0:4095];
  reg [31:0] pe56_lane18_strm1_tmp     ;
  reg [31:0] pe56_lane19_strm0 [0:4095];
  reg [31:0] pe56_lane19_strm0_tmp     ;
  reg [31:0] pe56_lane19_strm1 [0:4095];
  reg [31:0] pe56_lane19_strm1_tmp     ;
  reg [31:0] pe56_lane20_strm0 [0:4095];
  reg [31:0] pe56_lane20_strm0_tmp     ;
  reg [31:0] pe56_lane20_strm1 [0:4095];
  reg [31:0] pe56_lane20_strm1_tmp     ;
  reg [31:0] pe56_lane21_strm0 [0:4095];
  reg [31:0] pe56_lane21_strm0_tmp     ;
  reg [31:0] pe56_lane21_strm1 [0:4095];
  reg [31:0] pe56_lane21_strm1_tmp     ;
  reg [31:0] pe56_lane22_strm0 [0:4095];
  reg [31:0] pe56_lane22_strm0_tmp     ;
  reg [31:0] pe56_lane22_strm1 [0:4095];
  reg [31:0] pe56_lane22_strm1_tmp     ;
  reg [31:0] pe56_lane23_strm0 [0:4095];
  reg [31:0] pe56_lane23_strm0_tmp     ;
  reg [31:0] pe56_lane23_strm1 [0:4095];
  reg [31:0] pe56_lane23_strm1_tmp     ;
  reg [31:0] pe56_lane24_strm0 [0:4095];
  reg [31:0] pe56_lane24_strm0_tmp     ;
  reg [31:0] pe56_lane24_strm1 [0:4095];
  reg [31:0] pe56_lane24_strm1_tmp     ;
  reg [31:0] pe56_lane25_strm0 [0:4095];
  reg [31:0] pe56_lane25_strm0_tmp     ;
  reg [31:0] pe56_lane25_strm1 [0:4095];
  reg [31:0] pe56_lane25_strm1_tmp     ;
  reg [31:0] pe56_lane26_strm0 [0:4095];
  reg [31:0] pe56_lane26_strm0_tmp     ;
  reg [31:0] pe56_lane26_strm1 [0:4095];
  reg [31:0] pe56_lane26_strm1_tmp     ;
  reg [31:0] pe56_lane27_strm0 [0:4095];
  reg [31:0] pe56_lane27_strm0_tmp     ;
  reg [31:0] pe56_lane27_strm1 [0:4095];
  reg [31:0] pe56_lane27_strm1_tmp     ;
  reg [31:0] pe56_lane28_strm0 [0:4095];
  reg [31:0] pe56_lane28_strm0_tmp     ;
  reg [31:0] pe56_lane28_strm1 [0:4095];
  reg [31:0] pe56_lane28_strm1_tmp     ;
  reg [31:0] pe56_lane29_strm0 [0:4095];
  reg [31:0] pe56_lane29_strm0_tmp     ;
  reg [31:0] pe56_lane29_strm1 [0:4095];
  reg [31:0] pe56_lane29_strm1_tmp     ;
  reg [31:0] pe56_lane30_strm0 [0:4095];
  reg [31:0] pe56_lane30_strm0_tmp     ;
  reg [31:0] pe56_lane30_strm1 [0:4095];
  reg [31:0] pe56_lane30_strm1_tmp     ;
  reg [31:0] pe56_lane31_strm0 [0:4095];
  reg [31:0] pe56_lane31_strm0_tmp     ;
  reg [31:0] pe56_lane31_strm1 [0:4095];
  reg [31:0] pe56_lane31_strm1_tmp     ;
  reg [31:0] pe57_lane0_strm0 [0:4095];
  reg [31:0] pe57_lane0_strm0_tmp     ;
  reg [31:0] pe57_lane0_strm1 [0:4095];
  reg [31:0] pe57_lane0_strm1_tmp     ;
  reg [31:0] pe57_lane1_strm0 [0:4095];
  reg [31:0] pe57_lane1_strm0_tmp     ;
  reg [31:0] pe57_lane1_strm1 [0:4095];
  reg [31:0] pe57_lane1_strm1_tmp     ;
  reg [31:0] pe57_lane2_strm0 [0:4095];
  reg [31:0] pe57_lane2_strm0_tmp     ;
  reg [31:0] pe57_lane2_strm1 [0:4095];
  reg [31:0] pe57_lane2_strm1_tmp     ;
  reg [31:0] pe57_lane3_strm0 [0:4095];
  reg [31:0] pe57_lane3_strm0_tmp     ;
  reg [31:0] pe57_lane3_strm1 [0:4095];
  reg [31:0] pe57_lane3_strm1_tmp     ;
  reg [31:0] pe57_lane4_strm0 [0:4095];
  reg [31:0] pe57_lane4_strm0_tmp     ;
  reg [31:0] pe57_lane4_strm1 [0:4095];
  reg [31:0] pe57_lane4_strm1_tmp     ;
  reg [31:0] pe57_lane5_strm0 [0:4095];
  reg [31:0] pe57_lane5_strm0_tmp     ;
  reg [31:0] pe57_lane5_strm1 [0:4095];
  reg [31:0] pe57_lane5_strm1_tmp     ;
  reg [31:0] pe57_lane6_strm0 [0:4095];
  reg [31:0] pe57_lane6_strm0_tmp     ;
  reg [31:0] pe57_lane6_strm1 [0:4095];
  reg [31:0] pe57_lane6_strm1_tmp     ;
  reg [31:0] pe57_lane7_strm0 [0:4095];
  reg [31:0] pe57_lane7_strm0_tmp     ;
  reg [31:0] pe57_lane7_strm1 [0:4095];
  reg [31:0] pe57_lane7_strm1_tmp     ;
  reg [31:0] pe57_lane8_strm0 [0:4095];
  reg [31:0] pe57_lane8_strm0_tmp     ;
  reg [31:0] pe57_lane8_strm1 [0:4095];
  reg [31:0] pe57_lane8_strm1_tmp     ;
  reg [31:0] pe57_lane9_strm0 [0:4095];
  reg [31:0] pe57_lane9_strm0_tmp     ;
  reg [31:0] pe57_lane9_strm1 [0:4095];
  reg [31:0] pe57_lane9_strm1_tmp     ;
  reg [31:0] pe57_lane10_strm0 [0:4095];
  reg [31:0] pe57_lane10_strm0_tmp     ;
  reg [31:0] pe57_lane10_strm1 [0:4095];
  reg [31:0] pe57_lane10_strm1_tmp     ;
  reg [31:0] pe57_lane11_strm0 [0:4095];
  reg [31:0] pe57_lane11_strm0_tmp     ;
  reg [31:0] pe57_lane11_strm1 [0:4095];
  reg [31:0] pe57_lane11_strm1_tmp     ;
  reg [31:0] pe57_lane12_strm0 [0:4095];
  reg [31:0] pe57_lane12_strm0_tmp     ;
  reg [31:0] pe57_lane12_strm1 [0:4095];
  reg [31:0] pe57_lane12_strm1_tmp     ;
  reg [31:0] pe57_lane13_strm0 [0:4095];
  reg [31:0] pe57_lane13_strm0_tmp     ;
  reg [31:0] pe57_lane13_strm1 [0:4095];
  reg [31:0] pe57_lane13_strm1_tmp     ;
  reg [31:0] pe57_lane14_strm0 [0:4095];
  reg [31:0] pe57_lane14_strm0_tmp     ;
  reg [31:0] pe57_lane14_strm1 [0:4095];
  reg [31:0] pe57_lane14_strm1_tmp     ;
  reg [31:0] pe57_lane15_strm0 [0:4095];
  reg [31:0] pe57_lane15_strm0_tmp     ;
  reg [31:0] pe57_lane15_strm1 [0:4095];
  reg [31:0] pe57_lane15_strm1_tmp     ;
  reg [31:0] pe57_lane16_strm0 [0:4095];
  reg [31:0] pe57_lane16_strm0_tmp     ;
  reg [31:0] pe57_lane16_strm1 [0:4095];
  reg [31:0] pe57_lane16_strm1_tmp     ;
  reg [31:0] pe57_lane17_strm0 [0:4095];
  reg [31:0] pe57_lane17_strm0_tmp     ;
  reg [31:0] pe57_lane17_strm1 [0:4095];
  reg [31:0] pe57_lane17_strm1_tmp     ;
  reg [31:0] pe57_lane18_strm0 [0:4095];
  reg [31:0] pe57_lane18_strm0_tmp     ;
  reg [31:0] pe57_lane18_strm1 [0:4095];
  reg [31:0] pe57_lane18_strm1_tmp     ;
  reg [31:0] pe57_lane19_strm0 [0:4095];
  reg [31:0] pe57_lane19_strm0_tmp     ;
  reg [31:0] pe57_lane19_strm1 [0:4095];
  reg [31:0] pe57_lane19_strm1_tmp     ;
  reg [31:0] pe57_lane20_strm0 [0:4095];
  reg [31:0] pe57_lane20_strm0_tmp     ;
  reg [31:0] pe57_lane20_strm1 [0:4095];
  reg [31:0] pe57_lane20_strm1_tmp     ;
  reg [31:0] pe57_lane21_strm0 [0:4095];
  reg [31:0] pe57_lane21_strm0_tmp     ;
  reg [31:0] pe57_lane21_strm1 [0:4095];
  reg [31:0] pe57_lane21_strm1_tmp     ;
  reg [31:0] pe57_lane22_strm0 [0:4095];
  reg [31:0] pe57_lane22_strm0_tmp     ;
  reg [31:0] pe57_lane22_strm1 [0:4095];
  reg [31:0] pe57_lane22_strm1_tmp     ;
  reg [31:0] pe57_lane23_strm0 [0:4095];
  reg [31:0] pe57_lane23_strm0_tmp     ;
  reg [31:0] pe57_lane23_strm1 [0:4095];
  reg [31:0] pe57_lane23_strm1_tmp     ;
  reg [31:0] pe57_lane24_strm0 [0:4095];
  reg [31:0] pe57_lane24_strm0_tmp     ;
  reg [31:0] pe57_lane24_strm1 [0:4095];
  reg [31:0] pe57_lane24_strm1_tmp     ;
  reg [31:0] pe57_lane25_strm0 [0:4095];
  reg [31:0] pe57_lane25_strm0_tmp     ;
  reg [31:0] pe57_lane25_strm1 [0:4095];
  reg [31:0] pe57_lane25_strm1_tmp     ;
  reg [31:0] pe57_lane26_strm0 [0:4095];
  reg [31:0] pe57_lane26_strm0_tmp     ;
  reg [31:0] pe57_lane26_strm1 [0:4095];
  reg [31:0] pe57_lane26_strm1_tmp     ;
  reg [31:0] pe57_lane27_strm0 [0:4095];
  reg [31:0] pe57_lane27_strm0_tmp     ;
  reg [31:0] pe57_lane27_strm1 [0:4095];
  reg [31:0] pe57_lane27_strm1_tmp     ;
  reg [31:0] pe57_lane28_strm0 [0:4095];
  reg [31:0] pe57_lane28_strm0_tmp     ;
  reg [31:0] pe57_lane28_strm1 [0:4095];
  reg [31:0] pe57_lane28_strm1_tmp     ;
  reg [31:0] pe57_lane29_strm0 [0:4095];
  reg [31:0] pe57_lane29_strm0_tmp     ;
  reg [31:0] pe57_lane29_strm1 [0:4095];
  reg [31:0] pe57_lane29_strm1_tmp     ;
  reg [31:0] pe57_lane30_strm0 [0:4095];
  reg [31:0] pe57_lane30_strm0_tmp     ;
  reg [31:0] pe57_lane30_strm1 [0:4095];
  reg [31:0] pe57_lane30_strm1_tmp     ;
  reg [31:0] pe57_lane31_strm0 [0:4095];
  reg [31:0] pe57_lane31_strm0_tmp     ;
  reg [31:0] pe57_lane31_strm1 [0:4095];
  reg [31:0] pe57_lane31_strm1_tmp     ;
  reg [31:0] pe58_lane0_strm0 [0:4095];
  reg [31:0] pe58_lane0_strm0_tmp     ;
  reg [31:0] pe58_lane0_strm1 [0:4095];
  reg [31:0] pe58_lane0_strm1_tmp     ;
  reg [31:0] pe58_lane1_strm0 [0:4095];
  reg [31:0] pe58_lane1_strm0_tmp     ;
  reg [31:0] pe58_lane1_strm1 [0:4095];
  reg [31:0] pe58_lane1_strm1_tmp     ;
  reg [31:0] pe58_lane2_strm0 [0:4095];
  reg [31:0] pe58_lane2_strm0_tmp     ;
  reg [31:0] pe58_lane2_strm1 [0:4095];
  reg [31:0] pe58_lane2_strm1_tmp     ;
  reg [31:0] pe58_lane3_strm0 [0:4095];
  reg [31:0] pe58_lane3_strm0_tmp     ;
  reg [31:0] pe58_lane3_strm1 [0:4095];
  reg [31:0] pe58_lane3_strm1_tmp     ;
  reg [31:0] pe58_lane4_strm0 [0:4095];
  reg [31:0] pe58_lane4_strm0_tmp     ;
  reg [31:0] pe58_lane4_strm1 [0:4095];
  reg [31:0] pe58_lane4_strm1_tmp     ;
  reg [31:0] pe58_lane5_strm0 [0:4095];
  reg [31:0] pe58_lane5_strm0_tmp     ;
  reg [31:0] pe58_lane5_strm1 [0:4095];
  reg [31:0] pe58_lane5_strm1_tmp     ;
  reg [31:0] pe58_lane6_strm0 [0:4095];
  reg [31:0] pe58_lane6_strm0_tmp     ;
  reg [31:0] pe58_lane6_strm1 [0:4095];
  reg [31:0] pe58_lane6_strm1_tmp     ;
  reg [31:0] pe58_lane7_strm0 [0:4095];
  reg [31:0] pe58_lane7_strm0_tmp     ;
  reg [31:0] pe58_lane7_strm1 [0:4095];
  reg [31:0] pe58_lane7_strm1_tmp     ;
  reg [31:0] pe58_lane8_strm0 [0:4095];
  reg [31:0] pe58_lane8_strm0_tmp     ;
  reg [31:0] pe58_lane8_strm1 [0:4095];
  reg [31:0] pe58_lane8_strm1_tmp     ;
  reg [31:0] pe58_lane9_strm0 [0:4095];
  reg [31:0] pe58_lane9_strm0_tmp     ;
  reg [31:0] pe58_lane9_strm1 [0:4095];
  reg [31:0] pe58_lane9_strm1_tmp     ;
  reg [31:0] pe58_lane10_strm0 [0:4095];
  reg [31:0] pe58_lane10_strm0_tmp     ;
  reg [31:0] pe58_lane10_strm1 [0:4095];
  reg [31:0] pe58_lane10_strm1_tmp     ;
  reg [31:0] pe58_lane11_strm0 [0:4095];
  reg [31:0] pe58_lane11_strm0_tmp     ;
  reg [31:0] pe58_lane11_strm1 [0:4095];
  reg [31:0] pe58_lane11_strm1_tmp     ;
  reg [31:0] pe58_lane12_strm0 [0:4095];
  reg [31:0] pe58_lane12_strm0_tmp     ;
  reg [31:0] pe58_lane12_strm1 [0:4095];
  reg [31:0] pe58_lane12_strm1_tmp     ;
  reg [31:0] pe58_lane13_strm0 [0:4095];
  reg [31:0] pe58_lane13_strm0_tmp     ;
  reg [31:0] pe58_lane13_strm1 [0:4095];
  reg [31:0] pe58_lane13_strm1_tmp     ;
  reg [31:0] pe58_lane14_strm0 [0:4095];
  reg [31:0] pe58_lane14_strm0_tmp     ;
  reg [31:0] pe58_lane14_strm1 [0:4095];
  reg [31:0] pe58_lane14_strm1_tmp     ;
  reg [31:0] pe58_lane15_strm0 [0:4095];
  reg [31:0] pe58_lane15_strm0_tmp     ;
  reg [31:0] pe58_lane15_strm1 [0:4095];
  reg [31:0] pe58_lane15_strm1_tmp     ;
  reg [31:0] pe58_lane16_strm0 [0:4095];
  reg [31:0] pe58_lane16_strm0_tmp     ;
  reg [31:0] pe58_lane16_strm1 [0:4095];
  reg [31:0] pe58_lane16_strm1_tmp     ;
  reg [31:0] pe58_lane17_strm0 [0:4095];
  reg [31:0] pe58_lane17_strm0_tmp     ;
  reg [31:0] pe58_lane17_strm1 [0:4095];
  reg [31:0] pe58_lane17_strm1_tmp     ;
  reg [31:0] pe58_lane18_strm0 [0:4095];
  reg [31:0] pe58_lane18_strm0_tmp     ;
  reg [31:0] pe58_lane18_strm1 [0:4095];
  reg [31:0] pe58_lane18_strm1_tmp     ;
  reg [31:0] pe58_lane19_strm0 [0:4095];
  reg [31:0] pe58_lane19_strm0_tmp     ;
  reg [31:0] pe58_lane19_strm1 [0:4095];
  reg [31:0] pe58_lane19_strm1_tmp     ;
  reg [31:0] pe58_lane20_strm0 [0:4095];
  reg [31:0] pe58_lane20_strm0_tmp     ;
  reg [31:0] pe58_lane20_strm1 [0:4095];
  reg [31:0] pe58_lane20_strm1_tmp     ;
  reg [31:0] pe58_lane21_strm0 [0:4095];
  reg [31:0] pe58_lane21_strm0_tmp     ;
  reg [31:0] pe58_lane21_strm1 [0:4095];
  reg [31:0] pe58_lane21_strm1_tmp     ;
  reg [31:0] pe58_lane22_strm0 [0:4095];
  reg [31:0] pe58_lane22_strm0_tmp     ;
  reg [31:0] pe58_lane22_strm1 [0:4095];
  reg [31:0] pe58_lane22_strm1_tmp     ;
  reg [31:0] pe58_lane23_strm0 [0:4095];
  reg [31:0] pe58_lane23_strm0_tmp     ;
  reg [31:0] pe58_lane23_strm1 [0:4095];
  reg [31:0] pe58_lane23_strm1_tmp     ;
  reg [31:0] pe58_lane24_strm0 [0:4095];
  reg [31:0] pe58_lane24_strm0_tmp     ;
  reg [31:0] pe58_lane24_strm1 [0:4095];
  reg [31:0] pe58_lane24_strm1_tmp     ;
  reg [31:0] pe58_lane25_strm0 [0:4095];
  reg [31:0] pe58_lane25_strm0_tmp     ;
  reg [31:0] pe58_lane25_strm1 [0:4095];
  reg [31:0] pe58_lane25_strm1_tmp     ;
  reg [31:0] pe58_lane26_strm0 [0:4095];
  reg [31:0] pe58_lane26_strm0_tmp     ;
  reg [31:0] pe58_lane26_strm1 [0:4095];
  reg [31:0] pe58_lane26_strm1_tmp     ;
  reg [31:0] pe58_lane27_strm0 [0:4095];
  reg [31:0] pe58_lane27_strm0_tmp     ;
  reg [31:0] pe58_lane27_strm1 [0:4095];
  reg [31:0] pe58_lane27_strm1_tmp     ;
  reg [31:0] pe58_lane28_strm0 [0:4095];
  reg [31:0] pe58_lane28_strm0_tmp     ;
  reg [31:0] pe58_lane28_strm1 [0:4095];
  reg [31:0] pe58_lane28_strm1_tmp     ;
  reg [31:0] pe58_lane29_strm0 [0:4095];
  reg [31:0] pe58_lane29_strm0_tmp     ;
  reg [31:0] pe58_lane29_strm1 [0:4095];
  reg [31:0] pe58_lane29_strm1_tmp     ;
  reg [31:0] pe58_lane30_strm0 [0:4095];
  reg [31:0] pe58_lane30_strm0_tmp     ;
  reg [31:0] pe58_lane30_strm1 [0:4095];
  reg [31:0] pe58_lane30_strm1_tmp     ;
  reg [31:0] pe58_lane31_strm0 [0:4095];
  reg [31:0] pe58_lane31_strm0_tmp     ;
  reg [31:0] pe58_lane31_strm1 [0:4095];
  reg [31:0] pe58_lane31_strm1_tmp     ;
  reg [31:0] pe59_lane0_strm0 [0:4095];
  reg [31:0] pe59_lane0_strm0_tmp     ;
  reg [31:0] pe59_lane0_strm1 [0:4095];
  reg [31:0] pe59_lane0_strm1_tmp     ;
  reg [31:0] pe59_lane1_strm0 [0:4095];
  reg [31:0] pe59_lane1_strm0_tmp     ;
  reg [31:0] pe59_lane1_strm1 [0:4095];
  reg [31:0] pe59_lane1_strm1_tmp     ;
  reg [31:0] pe59_lane2_strm0 [0:4095];
  reg [31:0] pe59_lane2_strm0_tmp     ;
  reg [31:0] pe59_lane2_strm1 [0:4095];
  reg [31:0] pe59_lane2_strm1_tmp     ;
  reg [31:0] pe59_lane3_strm0 [0:4095];
  reg [31:0] pe59_lane3_strm0_tmp     ;
  reg [31:0] pe59_lane3_strm1 [0:4095];
  reg [31:0] pe59_lane3_strm1_tmp     ;
  reg [31:0] pe59_lane4_strm0 [0:4095];
  reg [31:0] pe59_lane4_strm0_tmp     ;
  reg [31:0] pe59_lane4_strm1 [0:4095];
  reg [31:0] pe59_lane4_strm1_tmp     ;
  reg [31:0] pe59_lane5_strm0 [0:4095];
  reg [31:0] pe59_lane5_strm0_tmp     ;
  reg [31:0] pe59_lane5_strm1 [0:4095];
  reg [31:0] pe59_lane5_strm1_tmp     ;
  reg [31:0] pe59_lane6_strm0 [0:4095];
  reg [31:0] pe59_lane6_strm0_tmp     ;
  reg [31:0] pe59_lane6_strm1 [0:4095];
  reg [31:0] pe59_lane6_strm1_tmp     ;
  reg [31:0] pe59_lane7_strm0 [0:4095];
  reg [31:0] pe59_lane7_strm0_tmp     ;
  reg [31:0] pe59_lane7_strm1 [0:4095];
  reg [31:0] pe59_lane7_strm1_tmp     ;
  reg [31:0] pe59_lane8_strm0 [0:4095];
  reg [31:0] pe59_lane8_strm0_tmp     ;
  reg [31:0] pe59_lane8_strm1 [0:4095];
  reg [31:0] pe59_lane8_strm1_tmp     ;
  reg [31:0] pe59_lane9_strm0 [0:4095];
  reg [31:0] pe59_lane9_strm0_tmp     ;
  reg [31:0] pe59_lane9_strm1 [0:4095];
  reg [31:0] pe59_lane9_strm1_tmp     ;
  reg [31:0] pe59_lane10_strm0 [0:4095];
  reg [31:0] pe59_lane10_strm0_tmp     ;
  reg [31:0] pe59_lane10_strm1 [0:4095];
  reg [31:0] pe59_lane10_strm1_tmp     ;
  reg [31:0] pe59_lane11_strm0 [0:4095];
  reg [31:0] pe59_lane11_strm0_tmp     ;
  reg [31:0] pe59_lane11_strm1 [0:4095];
  reg [31:0] pe59_lane11_strm1_tmp     ;
  reg [31:0] pe59_lane12_strm0 [0:4095];
  reg [31:0] pe59_lane12_strm0_tmp     ;
  reg [31:0] pe59_lane12_strm1 [0:4095];
  reg [31:0] pe59_lane12_strm1_tmp     ;
  reg [31:0] pe59_lane13_strm0 [0:4095];
  reg [31:0] pe59_lane13_strm0_tmp     ;
  reg [31:0] pe59_lane13_strm1 [0:4095];
  reg [31:0] pe59_lane13_strm1_tmp     ;
  reg [31:0] pe59_lane14_strm0 [0:4095];
  reg [31:0] pe59_lane14_strm0_tmp     ;
  reg [31:0] pe59_lane14_strm1 [0:4095];
  reg [31:0] pe59_lane14_strm1_tmp     ;
  reg [31:0] pe59_lane15_strm0 [0:4095];
  reg [31:0] pe59_lane15_strm0_tmp     ;
  reg [31:0] pe59_lane15_strm1 [0:4095];
  reg [31:0] pe59_lane15_strm1_tmp     ;
  reg [31:0] pe59_lane16_strm0 [0:4095];
  reg [31:0] pe59_lane16_strm0_tmp     ;
  reg [31:0] pe59_lane16_strm1 [0:4095];
  reg [31:0] pe59_lane16_strm1_tmp     ;
  reg [31:0] pe59_lane17_strm0 [0:4095];
  reg [31:0] pe59_lane17_strm0_tmp     ;
  reg [31:0] pe59_lane17_strm1 [0:4095];
  reg [31:0] pe59_lane17_strm1_tmp     ;
  reg [31:0] pe59_lane18_strm0 [0:4095];
  reg [31:0] pe59_lane18_strm0_tmp     ;
  reg [31:0] pe59_lane18_strm1 [0:4095];
  reg [31:0] pe59_lane18_strm1_tmp     ;
  reg [31:0] pe59_lane19_strm0 [0:4095];
  reg [31:0] pe59_lane19_strm0_tmp     ;
  reg [31:0] pe59_lane19_strm1 [0:4095];
  reg [31:0] pe59_lane19_strm1_tmp     ;
  reg [31:0] pe59_lane20_strm0 [0:4095];
  reg [31:0] pe59_lane20_strm0_tmp     ;
  reg [31:0] pe59_lane20_strm1 [0:4095];
  reg [31:0] pe59_lane20_strm1_tmp     ;
  reg [31:0] pe59_lane21_strm0 [0:4095];
  reg [31:0] pe59_lane21_strm0_tmp     ;
  reg [31:0] pe59_lane21_strm1 [0:4095];
  reg [31:0] pe59_lane21_strm1_tmp     ;
  reg [31:0] pe59_lane22_strm0 [0:4095];
  reg [31:0] pe59_lane22_strm0_tmp     ;
  reg [31:0] pe59_lane22_strm1 [0:4095];
  reg [31:0] pe59_lane22_strm1_tmp     ;
  reg [31:0] pe59_lane23_strm0 [0:4095];
  reg [31:0] pe59_lane23_strm0_tmp     ;
  reg [31:0] pe59_lane23_strm1 [0:4095];
  reg [31:0] pe59_lane23_strm1_tmp     ;
  reg [31:0] pe59_lane24_strm0 [0:4095];
  reg [31:0] pe59_lane24_strm0_tmp     ;
  reg [31:0] pe59_lane24_strm1 [0:4095];
  reg [31:0] pe59_lane24_strm1_tmp     ;
  reg [31:0] pe59_lane25_strm0 [0:4095];
  reg [31:0] pe59_lane25_strm0_tmp     ;
  reg [31:0] pe59_lane25_strm1 [0:4095];
  reg [31:0] pe59_lane25_strm1_tmp     ;
  reg [31:0] pe59_lane26_strm0 [0:4095];
  reg [31:0] pe59_lane26_strm0_tmp     ;
  reg [31:0] pe59_lane26_strm1 [0:4095];
  reg [31:0] pe59_lane26_strm1_tmp     ;
  reg [31:0] pe59_lane27_strm0 [0:4095];
  reg [31:0] pe59_lane27_strm0_tmp     ;
  reg [31:0] pe59_lane27_strm1 [0:4095];
  reg [31:0] pe59_lane27_strm1_tmp     ;
  reg [31:0] pe59_lane28_strm0 [0:4095];
  reg [31:0] pe59_lane28_strm0_tmp     ;
  reg [31:0] pe59_lane28_strm1 [0:4095];
  reg [31:0] pe59_lane28_strm1_tmp     ;
  reg [31:0] pe59_lane29_strm0 [0:4095];
  reg [31:0] pe59_lane29_strm0_tmp     ;
  reg [31:0] pe59_lane29_strm1 [0:4095];
  reg [31:0] pe59_lane29_strm1_tmp     ;
  reg [31:0] pe59_lane30_strm0 [0:4095];
  reg [31:0] pe59_lane30_strm0_tmp     ;
  reg [31:0] pe59_lane30_strm1 [0:4095];
  reg [31:0] pe59_lane30_strm1_tmp     ;
  reg [31:0] pe59_lane31_strm0 [0:4095];
  reg [31:0] pe59_lane31_strm0_tmp     ;
  reg [31:0] pe59_lane31_strm1 [0:4095];
  reg [31:0] pe59_lane31_strm1_tmp     ;
  reg [31:0] pe60_lane0_strm0 [0:4095];
  reg [31:0] pe60_lane0_strm0_tmp     ;
  reg [31:0] pe60_lane0_strm1 [0:4095];
  reg [31:0] pe60_lane0_strm1_tmp     ;
  reg [31:0] pe60_lane1_strm0 [0:4095];
  reg [31:0] pe60_lane1_strm0_tmp     ;
  reg [31:0] pe60_lane1_strm1 [0:4095];
  reg [31:0] pe60_lane1_strm1_tmp     ;
  reg [31:0] pe60_lane2_strm0 [0:4095];
  reg [31:0] pe60_lane2_strm0_tmp     ;
  reg [31:0] pe60_lane2_strm1 [0:4095];
  reg [31:0] pe60_lane2_strm1_tmp     ;
  reg [31:0] pe60_lane3_strm0 [0:4095];
  reg [31:0] pe60_lane3_strm0_tmp     ;
  reg [31:0] pe60_lane3_strm1 [0:4095];
  reg [31:0] pe60_lane3_strm1_tmp     ;
  reg [31:0] pe60_lane4_strm0 [0:4095];
  reg [31:0] pe60_lane4_strm0_tmp     ;
  reg [31:0] pe60_lane4_strm1 [0:4095];
  reg [31:0] pe60_lane4_strm1_tmp     ;
  reg [31:0] pe60_lane5_strm0 [0:4095];
  reg [31:0] pe60_lane5_strm0_tmp     ;
  reg [31:0] pe60_lane5_strm1 [0:4095];
  reg [31:0] pe60_lane5_strm1_tmp     ;
  reg [31:0] pe60_lane6_strm0 [0:4095];
  reg [31:0] pe60_lane6_strm0_tmp     ;
  reg [31:0] pe60_lane6_strm1 [0:4095];
  reg [31:0] pe60_lane6_strm1_tmp     ;
  reg [31:0] pe60_lane7_strm0 [0:4095];
  reg [31:0] pe60_lane7_strm0_tmp     ;
  reg [31:0] pe60_lane7_strm1 [0:4095];
  reg [31:0] pe60_lane7_strm1_tmp     ;
  reg [31:0] pe60_lane8_strm0 [0:4095];
  reg [31:0] pe60_lane8_strm0_tmp     ;
  reg [31:0] pe60_lane8_strm1 [0:4095];
  reg [31:0] pe60_lane8_strm1_tmp     ;
  reg [31:0] pe60_lane9_strm0 [0:4095];
  reg [31:0] pe60_lane9_strm0_tmp     ;
  reg [31:0] pe60_lane9_strm1 [0:4095];
  reg [31:0] pe60_lane9_strm1_tmp     ;
  reg [31:0] pe60_lane10_strm0 [0:4095];
  reg [31:0] pe60_lane10_strm0_tmp     ;
  reg [31:0] pe60_lane10_strm1 [0:4095];
  reg [31:0] pe60_lane10_strm1_tmp     ;
  reg [31:0] pe60_lane11_strm0 [0:4095];
  reg [31:0] pe60_lane11_strm0_tmp     ;
  reg [31:0] pe60_lane11_strm1 [0:4095];
  reg [31:0] pe60_lane11_strm1_tmp     ;
  reg [31:0] pe60_lane12_strm0 [0:4095];
  reg [31:0] pe60_lane12_strm0_tmp     ;
  reg [31:0] pe60_lane12_strm1 [0:4095];
  reg [31:0] pe60_lane12_strm1_tmp     ;
  reg [31:0] pe60_lane13_strm0 [0:4095];
  reg [31:0] pe60_lane13_strm0_tmp     ;
  reg [31:0] pe60_lane13_strm1 [0:4095];
  reg [31:0] pe60_lane13_strm1_tmp     ;
  reg [31:0] pe60_lane14_strm0 [0:4095];
  reg [31:0] pe60_lane14_strm0_tmp     ;
  reg [31:0] pe60_lane14_strm1 [0:4095];
  reg [31:0] pe60_lane14_strm1_tmp     ;
  reg [31:0] pe60_lane15_strm0 [0:4095];
  reg [31:0] pe60_lane15_strm0_tmp     ;
  reg [31:0] pe60_lane15_strm1 [0:4095];
  reg [31:0] pe60_lane15_strm1_tmp     ;
  reg [31:0] pe60_lane16_strm0 [0:4095];
  reg [31:0] pe60_lane16_strm0_tmp     ;
  reg [31:0] pe60_lane16_strm1 [0:4095];
  reg [31:0] pe60_lane16_strm1_tmp     ;
  reg [31:0] pe60_lane17_strm0 [0:4095];
  reg [31:0] pe60_lane17_strm0_tmp     ;
  reg [31:0] pe60_lane17_strm1 [0:4095];
  reg [31:0] pe60_lane17_strm1_tmp     ;
  reg [31:0] pe60_lane18_strm0 [0:4095];
  reg [31:0] pe60_lane18_strm0_tmp     ;
  reg [31:0] pe60_lane18_strm1 [0:4095];
  reg [31:0] pe60_lane18_strm1_tmp     ;
  reg [31:0] pe60_lane19_strm0 [0:4095];
  reg [31:0] pe60_lane19_strm0_tmp     ;
  reg [31:0] pe60_lane19_strm1 [0:4095];
  reg [31:0] pe60_lane19_strm1_tmp     ;
  reg [31:0] pe60_lane20_strm0 [0:4095];
  reg [31:0] pe60_lane20_strm0_tmp     ;
  reg [31:0] pe60_lane20_strm1 [0:4095];
  reg [31:0] pe60_lane20_strm1_tmp     ;
  reg [31:0] pe60_lane21_strm0 [0:4095];
  reg [31:0] pe60_lane21_strm0_tmp     ;
  reg [31:0] pe60_lane21_strm1 [0:4095];
  reg [31:0] pe60_lane21_strm1_tmp     ;
  reg [31:0] pe60_lane22_strm0 [0:4095];
  reg [31:0] pe60_lane22_strm0_tmp     ;
  reg [31:0] pe60_lane22_strm1 [0:4095];
  reg [31:0] pe60_lane22_strm1_tmp     ;
  reg [31:0] pe60_lane23_strm0 [0:4095];
  reg [31:0] pe60_lane23_strm0_tmp     ;
  reg [31:0] pe60_lane23_strm1 [0:4095];
  reg [31:0] pe60_lane23_strm1_tmp     ;
  reg [31:0] pe60_lane24_strm0 [0:4095];
  reg [31:0] pe60_lane24_strm0_tmp     ;
  reg [31:0] pe60_lane24_strm1 [0:4095];
  reg [31:0] pe60_lane24_strm1_tmp     ;
  reg [31:0] pe60_lane25_strm0 [0:4095];
  reg [31:0] pe60_lane25_strm0_tmp     ;
  reg [31:0] pe60_lane25_strm1 [0:4095];
  reg [31:0] pe60_lane25_strm1_tmp     ;
  reg [31:0] pe60_lane26_strm0 [0:4095];
  reg [31:0] pe60_lane26_strm0_tmp     ;
  reg [31:0] pe60_lane26_strm1 [0:4095];
  reg [31:0] pe60_lane26_strm1_tmp     ;
  reg [31:0] pe60_lane27_strm0 [0:4095];
  reg [31:0] pe60_lane27_strm0_tmp     ;
  reg [31:0] pe60_lane27_strm1 [0:4095];
  reg [31:0] pe60_lane27_strm1_tmp     ;
  reg [31:0] pe60_lane28_strm0 [0:4095];
  reg [31:0] pe60_lane28_strm0_tmp     ;
  reg [31:0] pe60_lane28_strm1 [0:4095];
  reg [31:0] pe60_lane28_strm1_tmp     ;
  reg [31:0] pe60_lane29_strm0 [0:4095];
  reg [31:0] pe60_lane29_strm0_tmp     ;
  reg [31:0] pe60_lane29_strm1 [0:4095];
  reg [31:0] pe60_lane29_strm1_tmp     ;
  reg [31:0] pe60_lane30_strm0 [0:4095];
  reg [31:0] pe60_lane30_strm0_tmp     ;
  reg [31:0] pe60_lane30_strm1 [0:4095];
  reg [31:0] pe60_lane30_strm1_tmp     ;
  reg [31:0] pe60_lane31_strm0 [0:4095];
  reg [31:0] pe60_lane31_strm0_tmp     ;
  reg [31:0] pe60_lane31_strm1 [0:4095];
  reg [31:0] pe60_lane31_strm1_tmp     ;
  reg [31:0] pe61_lane0_strm0 [0:4095];
  reg [31:0] pe61_lane0_strm0_tmp     ;
  reg [31:0] pe61_lane0_strm1 [0:4095];
  reg [31:0] pe61_lane0_strm1_tmp     ;
  reg [31:0] pe61_lane1_strm0 [0:4095];
  reg [31:0] pe61_lane1_strm0_tmp     ;
  reg [31:0] pe61_lane1_strm1 [0:4095];
  reg [31:0] pe61_lane1_strm1_tmp     ;
  reg [31:0] pe61_lane2_strm0 [0:4095];
  reg [31:0] pe61_lane2_strm0_tmp     ;
  reg [31:0] pe61_lane2_strm1 [0:4095];
  reg [31:0] pe61_lane2_strm1_tmp     ;
  reg [31:0] pe61_lane3_strm0 [0:4095];
  reg [31:0] pe61_lane3_strm0_tmp     ;
  reg [31:0] pe61_lane3_strm1 [0:4095];
  reg [31:0] pe61_lane3_strm1_tmp     ;
  reg [31:0] pe61_lane4_strm0 [0:4095];
  reg [31:0] pe61_lane4_strm0_tmp     ;
  reg [31:0] pe61_lane4_strm1 [0:4095];
  reg [31:0] pe61_lane4_strm1_tmp     ;
  reg [31:0] pe61_lane5_strm0 [0:4095];
  reg [31:0] pe61_lane5_strm0_tmp     ;
  reg [31:0] pe61_lane5_strm1 [0:4095];
  reg [31:0] pe61_lane5_strm1_tmp     ;
  reg [31:0] pe61_lane6_strm0 [0:4095];
  reg [31:0] pe61_lane6_strm0_tmp     ;
  reg [31:0] pe61_lane6_strm1 [0:4095];
  reg [31:0] pe61_lane6_strm1_tmp     ;
  reg [31:0] pe61_lane7_strm0 [0:4095];
  reg [31:0] pe61_lane7_strm0_tmp     ;
  reg [31:0] pe61_lane7_strm1 [0:4095];
  reg [31:0] pe61_lane7_strm1_tmp     ;
  reg [31:0] pe61_lane8_strm0 [0:4095];
  reg [31:0] pe61_lane8_strm0_tmp     ;
  reg [31:0] pe61_lane8_strm1 [0:4095];
  reg [31:0] pe61_lane8_strm1_tmp     ;
  reg [31:0] pe61_lane9_strm0 [0:4095];
  reg [31:0] pe61_lane9_strm0_tmp     ;
  reg [31:0] pe61_lane9_strm1 [0:4095];
  reg [31:0] pe61_lane9_strm1_tmp     ;
  reg [31:0] pe61_lane10_strm0 [0:4095];
  reg [31:0] pe61_lane10_strm0_tmp     ;
  reg [31:0] pe61_lane10_strm1 [0:4095];
  reg [31:0] pe61_lane10_strm1_tmp     ;
  reg [31:0] pe61_lane11_strm0 [0:4095];
  reg [31:0] pe61_lane11_strm0_tmp     ;
  reg [31:0] pe61_lane11_strm1 [0:4095];
  reg [31:0] pe61_lane11_strm1_tmp     ;
  reg [31:0] pe61_lane12_strm0 [0:4095];
  reg [31:0] pe61_lane12_strm0_tmp     ;
  reg [31:0] pe61_lane12_strm1 [0:4095];
  reg [31:0] pe61_lane12_strm1_tmp     ;
  reg [31:0] pe61_lane13_strm0 [0:4095];
  reg [31:0] pe61_lane13_strm0_tmp     ;
  reg [31:0] pe61_lane13_strm1 [0:4095];
  reg [31:0] pe61_lane13_strm1_tmp     ;
  reg [31:0] pe61_lane14_strm0 [0:4095];
  reg [31:0] pe61_lane14_strm0_tmp     ;
  reg [31:0] pe61_lane14_strm1 [0:4095];
  reg [31:0] pe61_lane14_strm1_tmp     ;
  reg [31:0] pe61_lane15_strm0 [0:4095];
  reg [31:0] pe61_lane15_strm0_tmp     ;
  reg [31:0] pe61_lane15_strm1 [0:4095];
  reg [31:0] pe61_lane15_strm1_tmp     ;
  reg [31:0] pe61_lane16_strm0 [0:4095];
  reg [31:0] pe61_lane16_strm0_tmp     ;
  reg [31:0] pe61_lane16_strm1 [0:4095];
  reg [31:0] pe61_lane16_strm1_tmp     ;
  reg [31:0] pe61_lane17_strm0 [0:4095];
  reg [31:0] pe61_lane17_strm0_tmp     ;
  reg [31:0] pe61_lane17_strm1 [0:4095];
  reg [31:0] pe61_lane17_strm1_tmp     ;
  reg [31:0] pe61_lane18_strm0 [0:4095];
  reg [31:0] pe61_lane18_strm0_tmp     ;
  reg [31:0] pe61_lane18_strm1 [0:4095];
  reg [31:0] pe61_lane18_strm1_tmp     ;
  reg [31:0] pe61_lane19_strm0 [0:4095];
  reg [31:0] pe61_lane19_strm0_tmp     ;
  reg [31:0] pe61_lane19_strm1 [0:4095];
  reg [31:0] pe61_lane19_strm1_tmp     ;
  reg [31:0] pe61_lane20_strm0 [0:4095];
  reg [31:0] pe61_lane20_strm0_tmp     ;
  reg [31:0] pe61_lane20_strm1 [0:4095];
  reg [31:0] pe61_lane20_strm1_tmp     ;
  reg [31:0] pe61_lane21_strm0 [0:4095];
  reg [31:0] pe61_lane21_strm0_tmp     ;
  reg [31:0] pe61_lane21_strm1 [0:4095];
  reg [31:0] pe61_lane21_strm1_tmp     ;
  reg [31:0] pe61_lane22_strm0 [0:4095];
  reg [31:0] pe61_lane22_strm0_tmp     ;
  reg [31:0] pe61_lane22_strm1 [0:4095];
  reg [31:0] pe61_lane22_strm1_tmp     ;
  reg [31:0] pe61_lane23_strm0 [0:4095];
  reg [31:0] pe61_lane23_strm0_tmp     ;
  reg [31:0] pe61_lane23_strm1 [0:4095];
  reg [31:0] pe61_lane23_strm1_tmp     ;
  reg [31:0] pe61_lane24_strm0 [0:4095];
  reg [31:0] pe61_lane24_strm0_tmp     ;
  reg [31:0] pe61_lane24_strm1 [0:4095];
  reg [31:0] pe61_lane24_strm1_tmp     ;
  reg [31:0] pe61_lane25_strm0 [0:4095];
  reg [31:0] pe61_lane25_strm0_tmp     ;
  reg [31:0] pe61_lane25_strm1 [0:4095];
  reg [31:0] pe61_lane25_strm1_tmp     ;
  reg [31:0] pe61_lane26_strm0 [0:4095];
  reg [31:0] pe61_lane26_strm0_tmp     ;
  reg [31:0] pe61_lane26_strm1 [0:4095];
  reg [31:0] pe61_lane26_strm1_tmp     ;
  reg [31:0] pe61_lane27_strm0 [0:4095];
  reg [31:0] pe61_lane27_strm0_tmp     ;
  reg [31:0] pe61_lane27_strm1 [0:4095];
  reg [31:0] pe61_lane27_strm1_tmp     ;
  reg [31:0] pe61_lane28_strm0 [0:4095];
  reg [31:0] pe61_lane28_strm0_tmp     ;
  reg [31:0] pe61_lane28_strm1 [0:4095];
  reg [31:0] pe61_lane28_strm1_tmp     ;
  reg [31:0] pe61_lane29_strm0 [0:4095];
  reg [31:0] pe61_lane29_strm0_tmp     ;
  reg [31:0] pe61_lane29_strm1 [0:4095];
  reg [31:0] pe61_lane29_strm1_tmp     ;
  reg [31:0] pe61_lane30_strm0 [0:4095];
  reg [31:0] pe61_lane30_strm0_tmp     ;
  reg [31:0] pe61_lane30_strm1 [0:4095];
  reg [31:0] pe61_lane30_strm1_tmp     ;
  reg [31:0] pe61_lane31_strm0 [0:4095];
  reg [31:0] pe61_lane31_strm0_tmp     ;
  reg [31:0] pe61_lane31_strm1 [0:4095];
  reg [31:0] pe61_lane31_strm1_tmp     ;
  reg [31:0] pe62_lane0_strm0 [0:4095];
  reg [31:0] pe62_lane0_strm0_tmp     ;
  reg [31:0] pe62_lane0_strm1 [0:4095];
  reg [31:0] pe62_lane0_strm1_tmp     ;
  reg [31:0] pe62_lane1_strm0 [0:4095];
  reg [31:0] pe62_lane1_strm0_tmp     ;
  reg [31:0] pe62_lane1_strm1 [0:4095];
  reg [31:0] pe62_lane1_strm1_tmp     ;
  reg [31:0] pe62_lane2_strm0 [0:4095];
  reg [31:0] pe62_lane2_strm0_tmp     ;
  reg [31:0] pe62_lane2_strm1 [0:4095];
  reg [31:0] pe62_lane2_strm1_tmp     ;
  reg [31:0] pe62_lane3_strm0 [0:4095];
  reg [31:0] pe62_lane3_strm0_tmp     ;
  reg [31:0] pe62_lane3_strm1 [0:4095];
  reg [31:0] pe62_lane3_strm1_tmp     ;
  reg [31:0] pe62_lane4_strm0 [0:4095];
  reg [31:0] pe62_lane4_strm0_tmp     ;
  reg [31:0] pe62_lane4_strm1 [0:4095];
  reg [31:0] pe62_lane4_strm1_tmp     ;
  reg [31:0] pe62_lane5_strm0 [0:4095];
  reg [31:0] pe62_lane5_strm0_tmp     ;
  reg [31:0] pe62_lane5_strm1 [0:4095];
  reg [31:0] pe62_lane5_strm1_tmp     ;
  reg [31:0] pe62_lane6_strm0 [0:4095];
  reg [31:0] pe62_lane6_strm0_tmp     ;
  reg [31:0] pe62_lane6_strm1 [0:4095];
  reg [31:0] pe62_lane6_strm1_tmp     ;
  reg [31:0] pe62_lane7_strm0 [0:4095];
  reg [31:0] pe62_lane7_strm0_tmp     ;
  reg [31:0] pe62_lane7_strm1 [0:4095];
  reg [31:0] pe62_lane7_strm1_tmp     ;
  reg [31:0] pe62_lane8_strm0 [0:4095];
  reg [31:0] pe62_lane8_strm0_tmp     ;
  reg [31:0] pe62_lane8_strm1 [0:4095];
  reg [31:0] pe62_lane8_strm1_tmp     ;
  reg [31:0] pe62_lane9_strm0 [0:4095];
  reg [31:0] pe62_lane9_strm0_tmp     ;
  reg [31:0] pe62_lane9_strm1 [0:4095];
  reg [31:0] pe62_lane9_strm1_tmp     ;
  reg [31:0] pe62_lane10_strm0 [0:4095];
  reg [31:0] pe62_lane10_strm0_tmp     ;
  reg [31:0] pe62_lane10_strm1 [0:4095];
  reg [31:0] pe62_lane10_strm1_tmp     ;
  reg [31:0] pe62_lane11_strm0 [0:4095];
  reg [31:0] pe62_lane11_strm0_tmp     ;
  reg [31:0] pe62_lane11_strm1 [0:4095];
  reg [31:0] pe62_lane11_strm1_tmp     ;
  reg [31:0] pe62_lane12_strm0 [0:4095];
  reg [31:0] pe62_lane12_strm0_tmp     ;
  reg [31:0] pe62_lane12_strm1 [0:4095];
  reg [31:0] pe62_lane12_strm1_tmp     ;
  reg [31:0] pe62_lane13_strm0 [0:4095];
  reg [31:0] pe62_lane13_strm0_tmp     ;
  reg [31:0] pe62_lane13_strm1 [0:4095];
  reg [31:0] pe62_lane13_strm1_tmp     ;
  reg [31:0] pe62_lane14_strm0 [0:4095];
  reg [31:0] pe62_lane14_strm0_tmp     ;
  reg [31:0] pe62_lane14_strm1 [0:4095];
  reg [31:0] pe62_lane14_strm1_tmp     ;
  reg [31:0] pe62_lane15_strm0 [0:4095];
  reg [31:0] pe62_lane15_strm0_tmp     ;
  reg [31:0] pe62_lane15_strm1 [0:4095];
  reg [31:0] pe62_lane15_strm1_tmp     ;
  reg [31:0] pe62_lane16_strm0 [0:4095];
  reg [31:0] pe62_lane16_strm0_tmp     ;
  reg [31:0] pe62_lane16_strm1 [0:4095];
  reg [31:0] pe62_lane16_strm1_tmp     ;
  reg [31:0] pe62_lane17_strm0 [0:4095];
  reg [31:0] pe62_lane17_strm0_tmp     ;
  reg [31:0] pe62_lane17_strm1 [0:4095];
  reg [31:0] pe62_lane17_strm1_tmp     ;
  reg [31:0] pe62_lane18_strm0 [0:4095];
  reg [31:0] pe62_lane18_strm0_tmp     ;
  reg [31:0] pe62_lane18_strm1 [0:4095];
  reg [31:0] pe62_lane18_strm1_tmp     ;
  reg [31:0] pe62_lane19_strm0 [0:4095];
  reg [31:0] pe62_lane19_strm0_tmp     ;
  reg [31:0] pe62_lane19_strm1 [0:4095];
  reg [31:0] pe62_lane19_strm1_tmp     ;
  reg [31:0] pe62_lane20_strm0 [0:4095];
  reg [31:0] pe62_lane20_strm0_tmp     ;
  reg [31:0] pe62_lane20_strm1 [0:4095];
  reg [31:0] pe62_lane20_strm1_tmp     ;
  reg [31:0] pe62_lane21_strm0 [0:4095];
  reg [31:0] pe62_lane21_strm0_tmp     ;
  reg [31:0] pe62_lane21_strm1 [0:4095];
  reg [31:0] pe62_lane21_strm1_tmp     ;
  reg [31:0] pe62_lane22_strm0 [0:4095];
  reg [31:0] pe62_lane22_strm0_tmp     ;
  reg [31:0] pe62_lane22_strm1 [0:4095];
  reg [31:0] pe62_lane22_strm1_tmp     ;
  reg [31:0] pe62_lane23_strm0 [0:4095];
  reg [31:0] pe62_lane23_strm0_tmp     ;
  reg [31:0] pe62_lane23_strm1 [0:4095];
  reg [31:0] pe62_lane23_strm1_tmp     ;
  reg [31:0] pe62_lane24_strm0 [0:4095];
  reg [31:0] pe62_lane24_strm0_tmp     ;
  reg [31:0] pe62_lane24_strm1 [0:4095];
  reg [31:0] pe62_lane24_strm1_tmp     ;
  reg [31:0] pe62_lane25_strm0 [0:4095];
  reg [31:0] pe62_lane25_strm0_tmp     ;
  reg [31:0] pe62_lane25_strm1 [0:4095];
  reg [31:0] pe62_lane25_strm1_tmp     ;
  reg [31:0] pe62_lane26_strm0 [0:4095];
  reg [31:0] pe62_lane26_strm0_tmp     ;
  reg [31:0] pe62_lane26_strm1 [0:4095];
  reg [31:0] pe62_lane26_strm1_tmp     ;
  reg [31:0] pe62_lane27_strm0 [0:4095];
  reg [31:0] pe62_lane27_strm0_tmp     ;
  reg [31:0] pe62_lane27_strm1 [0:4095];
  reg [31:0] pe62_lane27_strm1_tmp     ;
  reg [31:0] pe62_lane28_strm0 [0:4095];
  reg [31:0] pe62_lane28_strm0_tmp     ;
  reg [31:0] pe62_lane28_strm1 [0:4095];
  reg [31:0] pe62_lane28_strm1_tmp     ;
  reg [31:0] pe62_lane29_strm0 [0:4095];
  reg [31:0] pe62_lane29_strm0_tmp     ;
  reg [31:0] pe62_lane29_strm1 [0:4095];
  reg [31:0] pe62_lane29_strm1_tmp     ;
  reg [31:0] pe62_lane30_strm0 [0:4095];
  reg [31:0] pe62_lane30_strm0_tmp     ;
  reg [31:0] pe62_lane30_strm1 [0:4095];
  reg [31:0] pe62_lane30_strm1_tmp     ;
  reg [31:0] pe62_lane31_strm0 [0:4095];
  reg [31:0] pe62_lane31_strm0_tmp     ;
  reg [31:0] pe62_lane31_strm1 [0:4095];
  reg [31:0] pe62_lane31_strm1_tmp     ;
  reg [31:0] pe63_lane0_strm0 [0:4095];
  reg [31:0] pe63_lane0_strm0_tmp     ;
  reg [31:0] pe63_lane0_strm1 [0:4095];
  reg [31:0] pe63_lane0_strm1_tmp     ;
  reg [31:0] pe63_lane1_strm0 [0:4095];
  reg [31:0] pe63_lane1_strm0_tmp     ;
  reg [31:0] pe63_lane1_strm1 [0:4095];
  reg [31:0] pe63_lane1_strm1_tmp     ;
  reg [31:0] pe63_lane2_strm0 [0:4095];
  reg [31:0] pe63_lane2_strm0_tmp     ;
  reg [31:0] pe63_lane2_strm1 [0:4095];
  reg [31:0] pe63_lane2_strm1_tmp     ;
  reg [31:0] pe63_lane3_strm0 [0:4095];
  reg [31:0] pe63_lane3_strm0_tmp     ;
  reg [31:0] pe63_lane3_strm1 [0:4095];
  reg [31:0] pe63_lane3_strm1_tmp     ;
  reg [31:0] pe63_lane4_strm0 [0:4095];
  reg [31:0] pe63_lane4_strm0_tmp     ;
  reg [31:0] pe63_lane4_strm1 [0:4095];
  reg [31:0] pe63_lane4_strm1_tmp     ;
  reg [31:0] pe63_lane5_strm0 [0:4095];
  reg [31:0] pe63_lane5_strm0_tmp     ;
  reg [31:0] pe63_lane5_strm1 [0:4095];
  reg [31:0] pe63_lane5_strm1_tmp     ;
  reg [31:0] pe63_lane6_strm0 [0:4095];
  reg [31:0] pe63_lane6_strm0_tmp     ;
  reg [31:0] pe63_lane6_strm1 [0:4095];
  reg [31:0] pe63_lane6_strm1_tmp     ;
  reg [31:0] pe63_lane7_strm0 [0:4095];
  reg [31:0] pe63_lane7_strm0_tmp     ;
  reg [31:0] pe63_lane7_strm1 [0:4095];
  reg [31:0] pe63_lane7_strm1_tmp     ;
  reg [31:0] pe63_lane8_strm0 [0:4095];
  reg [31:0] pe63_lane8_strm0_tmp     ;
  reg [31:0] pe63_lane8_strm1 [0:4095];
  reg [31:0] pe63_lane8_strm1_tmp     ;
  reg [31:0] pe63_lane9_strm0 [0:4095];
  reg [31:0] pe63_lane9_strm0_tmp     ;
  reg [31:0] pe63_lane9_strm1 [0:4095];
  reg [31:0] pe63_lane9_strm1_tmp     ;
  reg [31:0] pe63_lane10_strm0 [0:4095];
  reg [31:0] pe63_lane10_strm0_tmp     ;
  reg [31:0] pe63_lane10_strm1 [0:4095];
  reg [31:0] pe63_lane10_strm1_tmp     ;
  reg [31:0] pe63_lane11_strm0 [0:4095];
  reg [31:0] pe63_lane11_strm0_tmp     ;
  reg [31:0] pe63_lane11_strm1 [0:4095];
  reg [31:0] pe63_lane11_strm1_tmp     ;
  reg [31:0] pe63_lane12_strm0 [0:4095];
  reg [31:0] pe63_lane12_strm0_tmp     ;
  reg [31:0] pe63_lane12_strm1 [0:4095];
  reg [31:0] pe63_lane12_strm1_tmp     ;
  reg [31:0] pe63_lane13_strm0 [0:4095];
  reg [31:0] pe63_lane13_strm0_tmp     ;
  reg [31:0] pe63_lane13_strm1 [0:4095];
  reg [31:0] pe63_lane13_strm1_tmp     ;
  reg [31:0] pe63_lane14_strm0 [0:4095];
  reg [31:0] pe63_lane14_strm0_tmp     ;
  reg [31:0] pe63_lane14_strm1 [0:4095];
  reg [31:0] pe63_lane14_strm1_tmp     ;
  reg [31:0] pe63_lane15_strm0 [0:4095];
  reg [31:0] pe63_lane15_strm0_tmp     ;
  reg [31:0] pe63_lane15_strm1 [0:4095];
  reg [31:0] pe63_lane15_strm1_tmp     ;
  reg [31:0] pe63_lane16_strm0 [0:4095];
  reg [31:0] pe63_lane16_strm0_tmp     ;
  reg [31:0] pe63_lane16_strm1 [0:4095];
  reg [31:0] pe63_lane16_strm1_tmp     ;
  reg [31:0] pe63_lane17_strm0 [0:4095];
  reg [31:0] pe63_lane17_strm0_tmp     ;
  reg [31:0] pe63_lane17_strm1 [0:4095];
  reg [31:0] pe63_lane17_strm1_tmp     ;
  reg [31:0] pe63_lane18_strm0 [0:4095];
  reg [31:0] pe63_lane18_strm0_tmp     ;
  reg [31:0] pe63_lane18_strm1 [0:4095];
  reg [31:0] pe63_lane18_strm1_tmp     ;
  reg [31:0] pe63_lane19_strm0 [0:4095];
  reg [31:0] pe63_lane19_strm0_tmp     ;
  reg [31:0] pe63_lane19_strm1 [0:4095];
  reg [31:0] pe63_lane19_strm1_tmp     ;
  reg [31:0] pe63_lane20_strm0 [0:4095];
  reg [31:0] pe63_lane20_strm0_tmp     ;
  reg [31:0] pe63_lane20_strm1 [0:4095];
  reg [31:0] pe63_lane20_strm1_tmp     ;
  reg [31:0] pe63_lane21_strm0 [0:4095];
  reg [31:0] pe63_lane21_strm0_tmp     ;
  reg [31:0] pe63_lane21_strm1 [0:4095];
  reg [31:0] pe63_lane21_strm1_tmp     ;
  reg [31:0] pe63_lane22_strm0 [0:4095];
  reg [31:0] pe63_lane22_strm0_tmp     ;
  reg [31:0] pe63_lane22_strm1 [0:4095];
  reg [31:0] pe63_lane22_strm1_tmp     ;
  reg [31:0] pe63_lane23_strm0 [0:4095];
  reg [31:0] pe63_lane23_strm0_tmp     ;
  reg [31:0] pe63_lane23_strm1 [0:4095];
  reg [31:0] pe63_lane23_strm1_tmp     ;
  reg [31:0] pe63_lane24_strm0 [0:4095];
  reg [31:0] pe63_lane24_strm0_tmp     ;
  reg [31:0] pe63_lane24_strm1 [0:4095];
  reg [31:0] pe63_lane24_strm1_tmp     ;
  reg [31:0] pe63_lane25_strm0 [0:4095];
  reg [31:0] pe63_lane25_strm0_tmp     ;
  reg [31:0] pe63_lane25_strm1 [0:4095];
  reg [31:0] pe63_lane25_strm1_tmp     ;
  reg [31:0] pe63_lane26_strm0 [0:4095];
  reg [31:0] pe63_lane26_strm0_tmp     ;
  reg [31:0] pe63_lane26_strm1 [0:4095];
  reg [31:0] pe63_lane26_strm1_tmp     ;
  reg [31:0] pe63_lane27_strm0 [0:4095];
  reg [31:0] pe63_lane27_strm0_tmp     ;
  reg [31:0] pe63_lane27_strm1 [0:4095];
  reg [31:0] pe63_lane27_strm1_tmp     ;
  reg [31:0] pe63_lane28_strm0 [0:4095];
  reg [31:0] pe63_lane28_strm0_tmp     ;
  reg [31:0] pe63_lane28_strm1 [0:4095];
  reg [31:0] pe63_lane28_strm1_tmp     ;
  reg [31:0] pe63_lane29_strm0 [0:4095];
  reg [31:0] pe63_lane29_strm0_tmp     ;
  reg [31:0] pe63_lane29_strm1 [0:4095];
  reg [31:0] pe63_lane29_strm1_tmp     ;
  reg [31:0] pe63_lane30_strm0 [0:4095];
  reg [31:0] pe63_lane30_strm0_tmp     ;
  reg [31:0] pe63_lane30_strm1 [0:4095];
  reg [31:0] pe63_lane30_strm1_tmp     ;
  reg [31:0] pe63_lane31_strm0 [0:4095];
  reg [31:0] pe63_lane31_strm0_tmp     ;
  reg [31:0] pe63_lane31_strm1 [0:4095];
  reg [31:0] pe63_lane31_strm1_tmp     ;