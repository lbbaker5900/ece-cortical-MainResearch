
  // OOB controls how the lanes are interpreted                                  
 assign    std__pe0__oob_cntl    =    mgr0__std__oob_cntl            ;
 assign    std__pe0__oob_valid   =    mgr0__std__oob_valid           ;
 assign    std__mgr0__oob_ready  =    pe0__std__oob_ready            ;
 assign    std__pe0__oob_type    =    mgr0__std__oob_type            ;
 assign    std__pe0__oob_data    =    mgr0__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe1__oob_cntl    =    mgr1__std__oob_cntl            ;
 assign    std__pe1__oob_valid   =    mgr1__std__oob_valid           ;
 assign    std__mgr1__oob_ready  =    pe1__std__oob_ready            ;
 assign    std__pe1__oob_type    =    mgr1__std__oob_type            ;
 assign    std__pe1__oob_data    =    mgr1__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe2__oob_cntl    =    mgr2__std__oob_cntl            ;
 assign    std__pe2__oob_valid   =    mgr2__std__oob_valid           ;
 assign    std__mgr2__oob_ready  =    pe2__std__oob_ready            ;
 assign    std__pe2__oob_type    =    mgr2__std__oob_type            ;
 assign    std__pe2__oob_data    =    mgr2__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe3__oob_cntl    =    mgr3__std__oob_cntl            ;
 assign    std__pe3__oob_valid   =    mgr3__std__oob_valid           ;
 assign    std__mgr3__oob_ready  =    pe3__std__oob_ready            ;
 assign    std__pe3__oob_type    =    mgr3__std__oob_type            ;
 assign    std__pe3__oob_data    =    mgr3__std__oob_data            ;
