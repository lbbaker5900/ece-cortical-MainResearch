
    wire                                           pe0__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe0__stu__cntl           ;
    wire                                           stu__pe0__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe0__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe0__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe0__stu__oob_data       ;

    wire                                           pe1__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe1__stu__cntl           ;
    wire                                           stu__pe1__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe1__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe1__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe1__stu__oob_data       ;

    wire                                           pe2__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe2__stu__cntl           ;
    wire                                           stu__pe2__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe2__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe2__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe2__stu__oob_data       ;

    wire                                           pe3__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe3__stu__cntl           ;
    wire                                           stu__pe3__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe3__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe3__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe3__stu__oob_data       ;

    wire                                           pe4__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe4__stu__cntl           ;
    wire                                           stu__pe4__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe4__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe4__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe4__stu__oob_data       ;

    wire                                           pe5__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe5__stu__cntl           ;
    wire                                           stu__pe5__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe5__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe5__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe5__stu__oob_data       ;

    wire                                           pe6__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe6__stu__cntl           ;
    wire                                           stu__pe6__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe6__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe6__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe6__stu__oob_data       ;

    wire                                           pe7__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe7__stu__cntl           ;
    wire                                           stu__pe7__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe7__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe7__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe7__stu__oob_data       ;

    wire                                           pe8__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe8__stu__cntl           ;
    wire                                           stu__pe8__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe8__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe8__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe8__stu__oob_data       ;

    wire                                           pe9__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe9__stu__cntl           ;
    wire                                           stu__pe9__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe9__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe9__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe9__stu__oob_data       ;

    wire                                           pe10__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe10__stu__cntl           ;
    wire                                           stu__pe10__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe10__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe10__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe10__stu__oob_data       ;

    wire                                           pe11__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe11__stu__cntl           ;
    wire                                           stu__pe11__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe11__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe11__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe11__stu__oob_data       ;

    wire                                           pe12__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe12__stu__cntl           ;
    wire                                           stu__pe12__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe12__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe12__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe12__stu__oob_data       ;

    wire                                           pe13__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe13__stu__cntl           ;
    wire                                           stu__pe13__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe13__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe13__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe13__stu__oob_data       ;

    wire                                           pe14__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe14__stu__cntl           ;
    wire                                           stu__pe14__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe14__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe14__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe14__stu__oob_data       ;

    wire                                           pe15__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe15__stu__cntl           ;
    wire                                           stu__pe15__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe15__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe15__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe15__stu__oob_data       ;

    wire                                           pe16__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe16__stu__cntl           ;
    wire                                           stu__pe16__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe16__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe16__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe16__stu__oob_data       ;

    wire                                           pe17__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe17__stu__cntl           ;
    wire                                           stu__pe17__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe17__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe17__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe17__stu__oob_data       ;

    wire                                           pe18__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe18__stu__cntl           ;
    wire                                           stu__pe18__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe18__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe18__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe18__stu__oob_data       ;

    wire                                           pe19__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe19__stu__cntl           ;
    wire                                           stu__pe19__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe19__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe19__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe19__stu__oob_data       ;

    wire                                           pe20__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe20__stu__cntl           ;
    wire                                           stu__pe20__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe20__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe20__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe20__stu__oob_data       ;

    wire                                           pe21__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe21__stu__cntl           ;
    wire                                           stu__pe21__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe21__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe21__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe21__stu__oob_data       ;

    wire                                           pe22__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe22__stu__cntl           ;
    wire                                           stu__pe22__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe22__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe22__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe22__stu__oob_data       ;

    wire                                           pe23__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe23__stu__cntl           ;
    wire                                           stu__pe23__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe23__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe23__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe23__stu__oob_data       ;

    wire                                           pe24__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe24__stu__cntl           ;
    wire                                           stu__pe24__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe24__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe24__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe24__stu__oob_data       ;

    wire                                           pe25__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe25__stu__cntl           ;
    wire                                           stu__pe25__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe25__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe25__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe25__stu__oob_data       ;

    wire                                           pe26__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe26__stu__cntl           ;
    wire                                           stu__pe26__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe26__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe26__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe26__stu__oob_data       ;

    wire                                           pe27__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe27__stu__cntl           ;
    wire                                           stu__pe27__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe27__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe27__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe27__stu__oob_data       ;

    wire                                           pe28__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe28__stu__cntl           ;
    wire                                           stu__pe28__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe28__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe28__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe28__stu__oob_data       ;

    wire                                           pe29__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe29__stu__cntl           ;
    wire                                           stu__pe29__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe29__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe29__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe29__stu__oob_data       ;

    wire                                           pe30__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe30__stu__cntl           ;
    wire                                           stu__pe30__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe30__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe30__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe30__stu__oob_data       ;

    wire                                           pe31__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe31__stu__cntl           ;
    wire                                           stu__pe31__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe31__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe31__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe31__stu__oob_data       ;

    wire                                           pe32__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe32__stu__cntl           ;
    wire                                           stu__pe32__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe32__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe32__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe32__stu__oob_data       ;

    wire                                           pe33__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe33__stu__cntl           ;
    wire                                           stu__pe33__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe33__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe33__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe33__stu__oob_data       ;

    wire                                           pe34__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe34__stu__cntl           ;
    wire                                           stu__pe34__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe34__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe34__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe34__stu__oob_data       ;

    wire                                           pe35__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe35__stu__cntl           ;
    wire                                           stu__pe35__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe35__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe35__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe35__stu__oob_data       ;

    wire                                           pe36__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe36__stu__cntl           ;
    wire                                           stu__pe36__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe36__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe36__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe36__stu__oob_data       ;

    wire                                           pe37__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe37__stu__cntl           ;
    wire                                           stu__pe37__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe37__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe37__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe37__stu__oob_data       ;

    wire                                           pe38__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe38__stu__cntl           ;
    wire                                           stu__pe38__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe38__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe38__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe38__stu__oob_data       ;

    wire                                           pe39__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe39__stu__cntl           ;
    wire                                           stu__pe39__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe39__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe39__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe39__stu__oob_data       ;

    wire                                           pe40__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe40__stu__cntl           ;
    wire                                           stu__pe40__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe40__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe40__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe40__stu__oob_data       ;

    wire                                           pe41__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe41__stu__cntl           ;
    wire                                           stu__pe41__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe41__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe41__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe41__stu__oob_data       ;

    wire                                           pe42__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe42__stu__cntl           ;
    wire                                           stu__pe42__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe42__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe42__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe42__stu__oob_data       ;

    wire                                           pe43__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe43__stu__cntl           ;
    wire                                           stu__pe43__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe43__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe43__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe43__stu__oob_data       ;

    wire                                           pe44__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe44__stu__cntl           ;
    wire                                           stu__pe44__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe44__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe44__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe44__stu__oob_data       ;

    wire                                           pe45__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe45__stu__cntl           ;
    wire                                           stu__pe45__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe45__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe45__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe45__stu__oob_data       ;

    wire                                           pe46__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe46__stu__cntl           ;
    wire                                           stu__pe46__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe46__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe46__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe46__stu__oob_data       ;

    wire                                           pe47__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe47__stu__cntl           ;
    wire                                           stu__pe47__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe47__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe47__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe47__stu__oob_data       ;

    wire                                           pe48__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe48__stu__cntl           ;
    wire                                           stu__pe48__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe48__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe48__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe48__stu__oob_data       ;

    wire                                           pe49__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe49__stu__cntl           ;
    wire                                           stu__pe49__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe49__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe49__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe49__stu__oob_data       ;

    wire                                           pe50__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe50__stu__cntl           ;
    wire                                           stu__pe50__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe50__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe50__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe50__stu__oob_data       ;

    wire                                           pe51__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe51__stu__cntl           ;
    wire                                           stu__pe51__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe51__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe51__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe51__stu__oob_data       ;

    wire                                           pe52__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe52__stu__cntl           ;
    wire                                           stu__pe52__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe52__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe52__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe52__stu__oob_data       ;

    wire                                           pe53__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe53__stu__cntl           ;
    wire                                           stu__pe53__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe53__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe53__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe53__stu__oob_data       ;

    wire                                           pe54__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe54__stu__cntl           ;
    wire                                           stu__pe54__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe54__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe54__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe54__stu__oob_data       ;

    wire                                           pe55__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe55__stu__cntl           ;
    wire                                           stu__pe55__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe55__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe55__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe55__stu__oob_data       ;

    wire                                           pe56__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe56__stu__cntl           ;
    wire                                           stu__pe56__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe56__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe56__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe56__stu__oob_data       ;

    wire                                           pe57__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe57__stu__cntl           ;
    wire                                           stu__pe57__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe57__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe57__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe57__stu__oob_data       ;

    wire                                           pe58__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe58__stu__cntl           ;
    wire                                           stu__pe58__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe58__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe58__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe58__stu__oob_data       ;

    wire                                           pe59__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe59__stu__cntl           ;
    wire                                           stu__pe59__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe59__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe59__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe59__stu__oob_data       ;

    wire                                           pe60__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe60__stu__cntl           ;
    wire                                           stu__pe60__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe60__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe60__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe60__stu__oob_data       ;

    wire                                           pe61__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe61__stu__cntl           ;
    wire                                           stu__pe61__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe61__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe61__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe61__stu__oob_data       ;

    wire                                           pe62__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe62__stu__cntl           ;
    wire                                           stu__pe62__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe62__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe62__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe62__stu__oob_data       ;

    wire                                           pe63__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe63__stu__cntl           ;
    wire                                           stu__pe63__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe63__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe63__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe63__stu__oob_data       ;

