
       // Aggregate Control-Path (cp) to NoC 
      .noc__cntl__cp_ready          ( noc__cntl__cp_ready         ), 
      .cntl__noc__cp_cntl           ( cntl__noc__cp_cntl          ), 
      .cntl__noc__cp_type           ( cntl__noc__cp_type          ), 
      .cntl__noc__cp_data           ( cntl__noc__cp_data          ), 
      .cntl__noc__cp_laneId         ( cntl__noc__cp_laneId        ), 
      .cntl__noc__cp_strmId         ( cntl__noc__cp_strmId        ), 
      .cntl__noc__cp_valid          ( cntl__noc__cp_valid         ), 
       // Aggregate Data-Path (cp) from NoC 
      .cntl__noc__cp_ready          ( cntl__noc__cp_ready         ), 
      .noc__cntl__cp_cntl           ( noc__cntl__cp_cntl          ), 
      .noc__cntl__cp_type           ( noc__cntl__cp_type          ), 
      .noc__cntl__cp_data           ( noc__cntl__cp_data          ), 
      .noc__cntl__cp_peId           ( noc__cntl__cp_peId          ), 
      .noc__cntl__cp_laneId         ( noc__cntl__cp_laneId        ), 
      .noc__cntl__cp_strmId         ( noc__cntl__cp_strmId        ), 
      .noc__cntl__cp_valid          ( noc__cntl__cp_valid         ), 

       // Aggregate Data-Path (dp) to NoC 
      .noc__cntl__dp_ready          ( noc__cntl__dp_ready         ), 
      .cntl__noc__dp_cntl           ( cntl__noc__dp_cntl          ), 
      .cntl__noc__dp_type           ( cntl__noc__dp_type          ), 
      .cntl__noc__dp_peId           ( cntl__noc__dp_peId          ), 
      .cntl__noc__dp_laneId         ( cntl__noc__dp_laneId        ), 
      .cntl__noc__dp_strmId         ( cntl__noc__dp_strmId        ), 
      .cntl__noc__dp_data           ( cntl__noc__dp_data          ), 
      .cntl__noc__dp_valid          ( cntl__noc__dp_valid         ), 
       // Aggregate Data-Path (dp) from NoC 
      .cntl__noc__dp_ready          ( cntl__noc__dp_ready         ), 
      .noc__cntl__dp_cntl           ( noc__cntl__dp_cntl          ), 
      .noc__cntl__dp_type           ( noc__cntl__dp_type          ), 
      .noc__cntl__dp_laneId         ( noc__cntl__dp_laneId        ), 
      .noc__cntl__dp_strmId         ( noc__cntl__dp_strmId        ), 
      .noc__cntl__dp_data           ( noc__cntl__dp_data          ), 
      .noc__cntl__dp_valid          ( noc__cntl__dp_valid         ), 
