
  // Lane 0, Stream 0
  assign stOp__sti__lane0_strm0_ready             =  stOp_lane[0].stOp__sti__strm0_ready  ;
  assign stOp_lane[0].sti__stOp__strm0_cntl       =  sti__stOp__lane0_strm0_cntl          ;
  assign stOp_lane[0].sti__stOp__strm0_data       =  sti__stOp__lane0_strm0_data          ;
  assign stOp_lane[0].sti__stOp__strm0_data_valid =  sti__stOp__lane0_strm0_data_valid    ;
  // Lane 1, Stream 0
  assign stOp__sti__lane1_strm0_ready             =  stOp_lane[1].stOp__sti__strm0_ready  ;
  assign stOp_lane[1].sti__stOp__strm0_cntl       =  sti__stOp__lane1_strm0_cntl          ;
  assign stOp_lane[1].sti__stOp__strm0_data       =  sti__stOp__lane1_strm0_data          ;
  assign stOp_lane[1].sti__stOp__strm0_data_valid =  sti__stOp__lane1_strm0_data_valid    ;
  // Lane 2, Stream 0
  assign stOp__sti__lane2_strm0_ready             =  stOp_lane[2].stOp__sti__strm0_ready  ;
  assign stOp_lane[2].sti__stOp__strm0_cntl       =  sti__stOp__lane2_strm0_cntl          ;
  assign stOp_lane[2].sti__stOp__strm0_data       =  sti__stOp__lane2_strm0_data          ;
  assign stOp_lane[2].sti__stOp__strm0_data_valid =  sti__stOp__lane2_strm0_data_valid    ;
  // Lane 3, Stream 0
  assign stOp__sti__lane3_strm0_ready             =  stOp_lane[3].stOp__sti__strm0_ready  ;
  assign stOp_lane[3].sti__stOp__strm0_cntl       =  sti__stOp__lane3_strm0_cntl          ;
  assign stOp_lane[3].sti__stOp__strm0_data       =  sti__stOp__lane3_strm0_data          ;
  assign stOp_lane[3].sti__stOp__strm0_data_valid =  sti__stOp__lane3_strm0_data_valid    ;
  // Lane 4, Stream 0
  assign stOp__sti__lane4_strm0_ready             =  stOp_lane[4].stOp__sti__strm0_ready  ;
  assign stOp_lane[4].sti__stOp__strm0_cntl       =  sti__stOp__lane4_strm0_cntl          ;
  assign stOp_lane[4].sti__stOp__strm0_data       =  sti__stOp__lane4_strm0_data          ;
  assign stOp_lane[4].sti__stOp__strm0_data_valid =  sti__stOp__lane4_strm0_data_valid    ;
  // Lane 5, Stream 0
  assign stOp__sti__lane5_strm0_ready             =  stOp_lane[5].stOp__sti__strm0_ready  ;
  assign stOp_lane[5].sti__stOp__strm0_cntl       =  sti__stOp__lane5_strm0_cntl          ;
  assign stOp_lane[5].sti__stOp__strm0_data       =  sti__stOp__lane5_strm0_data          ;
  assign stOp_lane[5].sti__stOp__strm0_data_valid =  sti__stOp__lane5_strm0_data_valid    ;
  // Lane 6, Stream 0
  assign stOp__sti__lane6_strm0_ready             =  stOp_lane[6].stOp__sti__strm0_ready  ;
  assign stOp_lane[6].sti__stOp__strm0_cntl       =  sti__stOp__lane6_strm0_cntl          ;
  assign stOp_lane[6].sti__stOp__strm0_data       =  sti__stOp__lane6_strm0_data          ;
  assign stOp_lane[6].sti__stOp__strm0_data_valid =  sti__stOp__lane6_strm0_data_valid    ;
  // Lane 7, Stream 0
  assign stOp__sti__lane7_strm0_ready             =  stOp_lane[7].stOp__sti__strm0_ready  ;
  assign stOp_lane[7].sti__stOp__strm0_cntl       =  sti__stOp__lane7_strm0_cntl          ;
  assign stOp_lane[7].sti__stOp__strm0_data       =  sti__stOp__lane7_strm0_data          ;
  assign stOp_lane[7].sti__stOp__strm0_data_valid =  sti__stOp__lane7_strm0_data_valid    ;
  // Lane 8, Stream 0
  assign stOp__sti__lane8_strm0_ready             =  stOp_lane[8].stOp__sti__strm0_ready  ;
  assign stOp_lane[8].sti__stOp__strm0_cntl       =  sti__stOp__lane8_strm0_cntl          ;
  assign stOp_lane[8].sti__stOp__strm0_data       =  sti__stOp__lane8_strm0_data          ;
  assign stOp_lane[8].sti__stOp__strm0_data_valid =  sti__stOp__lane8_strm0_data_valid    ;
  // Lane 9, Stream 0
  assign stOp__sti__lane9_strm0_ready             =  stOp_lane[9].stOp__sti__strm0_ready  ;
  assign stOp_lane[9].sti__stOp__strm0_cntl       =  sti__stOp__lane9_strm0_cntl          ;
  assign stOp_lane[9].sti__stOp__strm0_data       =  sti__stOp__lane9_strm0_data          ;
  assign stOp_lane[9].sti__stOp__strm0_data_valid =  sti__stOp__lane9_strm0_data_valid    ;
  // Lane 10, Stream 0
  assign stOp__sti__lane10_strm0_ready             =  stOp_lane[10].stOp__sti__strm0_ready  ;
  assign stOp_lane[10].sti__stOp__strm0_cntl       =  sti__stOp__lane10_strm0_cntl          ;
  assign stOp_lane[10].sti__stOp__strm0_data       =  sti__stOp__lane10_strm0_data          ;
  assign stOp_lane[10].sti__stOp__strm0_data_valid =  sti__stOp__lane10_strm0_data_valid    ;
  // Lane 11, Stream 0
  assign stOp__sti__lane11_strm0_ready             =  stOp_lane[11].stOp__sti__strm0_ready  ;
  assign stOp_lane[11].sti__stOp__strm0_cntl       =  sti__stOp__lane11_strm0_cntl          ;
  assign stOp_lane[11].sti__stOp__strm0_data       =  sti__stOp__lane11_strm0_data          ;
  assign stOp_lane[11].sti__stOp__strm0_data_valid =  sti__stOp__lane11_strm0_data_valid    ;
  // Lane 12, Stream 0
  assign stOp__sti__lane12_strm0_ready             =  stOp_lane[12].stOp__sti__strm0_ready  ;
  assign stOp_lane[12].sti__stOp__strm0_cntl       =  sti__stOp__lane12_strm0_cntl          ;
  assign stOp_lane[12].sti__stOp__strm0_data       =  sti__stOp__lane12_strm0_data          ;
  assign stOp_lane[12].sti__stOp__strm0_data_valid =  sti__stOp__lane12_strm0_data_valid    ;
  // Lane 13, Stream 0
  assign stOp__sti__lane13_strm0_ready             =  stOp_lane[13].stOp__sti__strm0_ready  ;
  assign stOp_lane[13].sti__stOp__strm0_cntl       =  sti__stOp__lane13_strm0_cntl          ;
  assign stOp_lane[13].sti__stOp__strm0_data       =  sti__stOp__lane13_strm0_data          ;
  assign stOp_lane[13].sti__stOp__strm0_data_valid =  sti__stOp__lane13_strm0_data_valid    ;
  // Lane 14, Stream 0
  assign stOp__sti__lane14_strm0_ready             =  stOp_lane[14].stOp__sti__strm0_ready  ;
  assign stOp_lane[14].sti__stOp__strm0_cntl       =  sti__stOp__lane14_strm0_cntl          ;
  assign stOp_lane[14].sti__stOp__strm0_data       =  sti__stOp__lane14_strm0_data          ;
  assign stOp_lane[14].sti__stOp__strm0_data_valid =  sti__stOp__lane14_strm0_data_valid    ;
  // Lane 15, Stream 0
  assign stOp__sti__lane15_strm0_ready             =  stOp_lane[15].stOp__sti__strm0_ready  ;
  assign stOp_lane[15].sti__stOp__strm0_cntl       =  sti__stOp__lane15_strm0_cntl          ;
  assign stOp_lane[15].sti__stOp__strm0_data       =  sti__stOp__lane15_strm0_data          ;
  assign stOp_lane[15].sti__stOp__strm0_data_valid =  sti__stOp__lane15_strm0_data_valid    ;
  // Lane 16, Stream 0
  assign stOp__sti__lane16_strm0_ready             =  stOp_lane[16].stOp__sti__strm0_ready  ;
  assign stOp_lane[16].sti__stOp__strm0_cntl       =  sti__stOp__lane16_strm0_cntl          ;
  assign stOp_lane[16].sti__stOp__strm0_data       =  sti__stOp__lane16_strm0_data          ;
  assign stOp_lane[16].sti__stOp__strm0_data_valid =  sti__stOp__lane16_strm0_data_valid    ;
  // Lane 17, Stream 0
  assign stOp__sti__lane17_strm0_ready             =  stOp_lane[17].stOp__sti__strm0_ready  ;
  assign stOp_lane[17].sti__stOp__strm0_cntl       =  sti__stOp__lane17_strm0_cntl          ;
  assign stOp_lane[17].sti__stOp__strm0_data       =  sti__stOp__lane17_strm0_data          ;
  assign stOp_lane[17].sti__stOp__strm0_data_valid =  sti__stOp__lane17_strm0_data_valid    ;
  // Lane 18, Stream 0
  assign stOp__sti__lane18_strm0_ready             =  stOp_lane[18].stOp__sti__strm0_ready  ;
  assign stOp_lane[18].sti__stOp__strm0_cntl       =  sti__stOp__lane18_strm0_cntl          ;
  assign stOp_lane[18].sti__stOp__strm0_data       =  sti__stOp__lane18_strm0_data          ;
  assign stOp_lane[18].sti__stOp__strm0_data_valid =  sti__stOp__lane18_strm0_data_valid    ;
  // Lane 19, Stream 0
  assign stOp__sti__lane19_strm0_ready             =  stOp_lane[19].stOp__sti__strm0_ready  ;
  assign stOp_lane[19].sti__stOp__strm0_cntl       =  sti__stOp__lane19_strm0_cntl          ;
  assign stOp_lane[19].sti__stOp__strm0_data       =  sti__stOp__lane19_strm0_data          ;
  assign stOp_lane[19].sti__stOp__strm0_data_valid =  sti__stOp__lane19_strm0_data_valid    ;
  // Lane 20, Stream 0
  assign stOp__sti__lane20_strm0_ready             =  stOp_lane[20].stOp__sti__strm0_ready  ;
  assign stOp_lane[20].sti__stOp__strm0_cntl       =  sti__stOp__lane20_strm0_cntl          ;
  assign stOp_lane[20].sti__stOp__strm0_data       =  sti__stOp__lane20_strm0_data          ;
  assign stOp_lane[20].sti__stOp__strm0_data_valid =  sti__stOp__lane20_strm0_data_valid    ;
  // Lane 21, Stream 0
  assign stOp__sti__lane21_strm0_ready             =  stOp_lane[21].stOp__sti__strm0_ready  ;
  assign stOp_lane[21].sti__stOp__strm0_cntl       =  sti__stOp__lane21_strm0_cntl          ;
  assign stOp_lane[21].sti__stOp__strm0_data       =  sti__stOp__lane21_strm0_data          ;
  assign stOp_lane[21].sti__stOp__strm0_data_valid =  sti__stOp__lane21_strm0_data_valid    ;
  // Lane 22, Stream 0
  assign stOp__sti__lane22_strm0_ready             =  stOp_lane[22].stOp__sti__strm0_ready  ;
  assign stOp_lane[22].sti__stOp__strm0_cntl       =  sti__stOp__lane22_strm0_cntl          ;
  assign stOp_lane[22].sti__stOp__strm0_data       =  sti__stOp__lane22_strm0_data          ;
  assign stOp_lane[22].sti__stOp__strm0_data_valid =  sti__stOp__lane22_strm0_data_valid    ;
  // Lane 23, Stream 0
  assign stOp__sti__lane23_strm0_ready             =  stOp_lane[23].stOp__sti__strm0_ready  ;
  assign stOp_lane[23].sti__stOp__strm0_cntl       =  sti__stOp__lane23_strm0_cntl          ;
  assign stOp_lane[23].sti__stOp__strm0_data       =  sti__stOp__lane23_strm0_data          ;
  assign stOp_lane[23].sti__stOp__strm0_data_valid =  sti__stOp__lane23_strm0_data_valid    ;
  // Lane 24, Stream 0
  assign stOp__sti__lane24_strm0_ready             =  stOp_lane[24].stOp__sti__strm0_ready  ;
  assign stOp_lane[24].sti__stOp__strm0_cntl       =  sti__stOp__lane24_strm0_cntl          ;
  assign stOp_lane[24].sti__stOp__strm0_data       =  sti__stOp__lane24_strm0_data          ;
  assign stOp_lane[24].sti__stOp__strm0_data_valid =  sti__stOp__lane24_strm0_data_valid    ;
  // Lane 25, Stream 0
  assign stOp__sti__lane25_strm0_ready             =  stOp_lane[25].stOp__sti__strm0_ready  ;
  assign stOp_lane[25].sti__stOp__strm0_cntl       =  sti__stOp__lane25_strm0_cntl          ;
  assign stOp_lane[25].sti__stOp__strm0_data       =  sti__stOp__lane25_strm0_data          ;
  assign stOp_lane[25].sti__stOp__strm0_data_valid =  sti__stOp__lane25_strm0_data_valid    ;
  // Lane 26, Stream 0
  assign stOp__sti__lane26_strm0_ready             =  stOp_lane[26].stOp__sti__strm0_ready  ;
  assign stOp_lane[26].sti__stOp__strm0_cntl       =  sti__stOp__lane26_strm0_cntl          ;
  assign stOp_lane[26].sti__stOp__strm0_data       =  sti__stOp__lane26_strm0_data          ;
  assign stOp_lane[26].sti__stOp__strm0_data_valid =  sti__stOp__lane26_strm0_data_valid    ;
  // Lane 27, Stream 0
  assign stOp__sti__lane27_strm0_ready             =  stOp_lane[27].stOp__sti__strm0_ready  ;
  assign stOp_lane[27].sti__stOp__strm0_cntl       =  sti__stOp__lane27_strm0_cntl          ;
  assign stOp_lane[27].sti__stOp__strm0_data       =  sti__stOp__lane27_strm0_data          ;
  assign stOp_lane[27].sti__stOp__strm0_data_valid =  sti__stOp__lane27_strm0_data_valid    ;
  // Lane 28, Stream 0
  assign stOp__sti__lane28_strm0_ready             =  stOp_lane[28].stOp__sti__strm0_ready  ;
  assign stOp_lane[28].sti__stOp__strm0_cntl       =  sti__stOp__lane28_strm0_cntl          ;
  assign stOp_lane[28].sti__stOp__strm0_data       =  sti__stOp__lane28_strm0_data          ;
  assign stOp_lane[28].sti__stOp__strm0_data_valid =  sti__stOp__lane28_strm0_data_valid    ;
  // Lane 29, Stream 0
  assign stOp__sti__lane29_strm0_ready             =  stOp_lane[29].stOp__sti__strm0_ready  ;
  assign stOp_lane[29].sti__stOp__strm0_cntl       =  sti__stOp__lane29_strm0_cntl          ;
  assign stOp_lane[29].sti__stOp__strm0_data       =  sti__stOp__lane29_strm0_data          ;
  assign stOp_lane[29].sti__stOp__strm0_data_valid =  sti__stOp__lane29_strm0_data_valid    ;
  // Lane 30, Stream 0
  assign stOp__sti__lane30_strm0_ready             =  stOp_lane[30].stOp__sti__strm0_ready  ;
  assign stOp_lane[30].sti__stOp__strm0_cntl       =  sti__stOp__lane30_strm0_cntl          ;
  assign stOp_lane[30].sti__stOp__strm0_data       =  sti__stOp__lane30_strm0_data          ;
  assign stOp_lane[30].sti__stOp__strm0_data_valid =  sti__stOp__lane30_strm0_data_valid    ;
  // Lane 31, Stream 0
  assign stOp__sti__lane31_strm0_ready             =  stOp_lane[31].stOp__sti__strm0_ready  ;
  assign stOp_lane[31].sti__stOp__strm0_cntl       =  sti__stOp__lane31_strm0_cntl          ;
  assign stOp_lane[31].sti__stOp__strm0_data       =  sti__stOp__lane31_strm0_data          ;
  assign stOp_lane[31].sti__stOp__strm0_data_valid =  sti__stOp__lane31_strm0_data_valid    ;

  // Lane 0, Stream 1
  assign stOp__sti__lane0_strm1_ready             =  stOp_lane[0].stOp__sti__strm1_ready  ;
  assign stOp_lane[0].sti__stOp__strm1_cntl       =  sti__stOp__lane0_strm1_cntl          ;
  assign stOp_lane[0].sti__stOp__strm1_data       =  sti__stOp__lane0_strm1_data          ;
  assign stOp_lane[0].sti__stOp__strm1_data_valid =  sti__stOp__lane0_strm1_data_valid    ;
  // Lane 1, Stream 1
  assign stOp__sti__lane1_strm1_ready             =  stOp_lane[1].stOp__sti__strm1_ready  ;
  assign stOp_lane[1].sti__stOp__strm1_cntl       =  sti__stOp__lane1_strm1_cntl          ;
  assign stOp_lane[1].sti__stOp__strm1_data       =  sti__stOp__lane1_strm1_data          ;
  assign stOp_lane[1].sti__stOp__strm1_data_valid =  sti__stOp__lane1_strm1_data_valid    ;
  // Lane 2, Stream 1
  assign stOp__sti__lane2_strm1_ready             =  stOp_lane[2].stOp__sti__strm1_ready  ;
  assign stOp_lane[2].sti__stOp__strm1_cntl       =  sti__stOp__lane2_strm1_cntl          ;
  assign stOp_lane[2].sti__stOp__strm1_data       =  sti__stOp__lane2_strm1_data          ;
  assign stOp_lane[2].sti__stOp__strm1_data_valid =  sti__stOp__lane2_strm1_data_valid    ;
  // Lane 3, Stream 1
  assign stOp__sti__lane3_strm1_ready             =  stOp_lane[3].stOp__sti__strm1_ready  ;
  assign stOp_lane[3].sti__stOp__strm1_cntl       =  sti__stOp__lane3_strm1_cntl          ;
  assign stOp_lane[3].sti__stOp__strm1_data       =  sti__stOp__lane3_strm1_data          ;
  assign stOp_lane[3].sti__stOp__strm1_data_valid =  sti__stOp__lane3_strm1_data_valid    ;
  // Lane 4, Stream 1
  assign stOp__sti__lane4_strm1_ready             =  stOp_lane[4].stOp__sti__strm1_ready  ;
  assign stOp_lane[4].sti__stOp__strm1_cntl       =  sti__stOp__lane4_strm1_cntl          ;
  assign stOp_lane[4].sti__stOp__strm1_data       =  sti__stOp__lane4_strm1_data          ;
  assign stOp_lane[4].sti__stOp__strm1_data_valid =  sti__stOp__lane4_strm1_data_valid    ;
  // Lane 5, Stream 1
  assign stOp__sti__lane5_strm1_ready             =  stOp_lane[5].stOp__sti__strm1_ready  ;
  assign stOp_lane[5].sti__stOp__strm1_cntl       =  sti__stOp__lane5_strm1_cntl          ;
  assign stOp_lane[5].sti__stOp__strm1_data       =  sti__stOp__lane5_strm1_data          ;
  assign stOp_lane[5].sti__stOp__strm1_data_valid =  sti__stOp__lane5_strm1_data_valid    ;
  // Lane 6, Stream 1
  assign stOp__sti__lane6_strm1_ready             =  stOp_lane[6].stOp__sti__strm1_ready  ;
  assign stOp_lane[6].sti__stOp__strm1_cntl       =  sti__stOp__lane6_strm1_cntl          ;
  assign stOp_lane[6].sti__stOp__strm1_data       =  sti__stOp__lane6_strm1_data          ;
  assign stOp_lane[6].sti__stOp__strm1_data_valid =  sti__stOp__lane6_strm1_data_valid    ;
  // Lane 7, Stream 1
  assign stOp__sti__lane7_strm1_ready             =  stOp_lane[7].stOp__sti__strm1_ready  ;
  assign stOp_lane[7].sti__stOp__strm1_cntl       =  sti__stOp__lane7_strm1_cntl          ;
  assign stOp_lane[7].sti__stOp__strm1_data       =  sti__stOp__lane7_strm1_data          ;
  assign stOp_lane[7].sti__stOp__strm1_data_valid =  sti__stOp__lane7_strm1_data_valid    ;
  // Lane 8, Stream 1
  assign stOp__sti__lane8_strm1_ready             =  stOp_lane[8].stOp__sti__strm1_ready  ;
  assign stOp_lane[8].sti__stOp__strm1_cntl       =  sti__stOp__lane8_strm1_cntl          ;
  assign stOp_lane[8].sti__stOp__strm1_data       =  sti__stOp__lane8_strm1_data          ;
  assign stOp_lane[8].sti__stOp__strm1_data_valid =  sti__stOp__lane8_strm1_data_valid    ;
  // Lane 9, Stream 1
  assign stOp__sti__lane9_strm1_ready             =  stOp_lane[9].stOp__sti__strm1_ready  ;
  assign stOp_lane[9].sti__stOp__strm1_cntl       =  sti__stOp__lane9_strm1_cntl          ;
  assign stOp_lane[9].sti__stOp__strm1_data       =  sti__stOp__lane9_strm1_data          ;
  assign stOp_lane[9].sti__stOp__strm1_data_valid =  sti__stOp__lane9_strm1_data_valid    ;
  // Lane 10, Stream 1
  assign stOp__sti__lane10_strm1_ready             =  stOp_lane[10].stOp__sti__strm1_ready  ;
  assign stOp_lane[10].sti__stOp__strm1_cntl       =  sti__stOp__lane10_strm1_cntl          ;
  assign stOp_lane[10].sti__stOp__strm1_data       =  sti__stOp__lane10_strm1_data          ;
  assign stOp_lane[10].sti__stOp__strm1_data_valid =  sti__stOp__lane10_strm1_data_valid    ;
  // Lane 11, Stream 1
  assign stOp__sti__lane11_strm1_ready             =  stOp_lane[11].stOp__sti__strm1_ready  ;
  assign stOp_lane[11].sti__stOp__strm1_cntl       =  sti__stOp__lane11_strm1_cntl          ;
  assign stOp_lane[11].sti__stOp__strm1_data       =  sti__stOp__lane11_strm1_data          ;
  assign stOp_lane[11].sti__stOp__strm1_data_valid =  sti__stOp__lane11_strm1_data_valid    ;
  // Lane 12, Stream 1
  assign stOp__sti__lane12_strm1_ready             =  stOp_lane[12].stOp__sti__strm1_ready  ;
  assign stOp_lane[12].sti__stOp__strm1_cntl       =  sti__stOp__lane12_strm1_cntl          ;
  assign stOp_lane[12].sti__stOp__strm1_data       =  sti__stOp__lane12_strm1_data          ;
  assign stOp_lane[12].sti__stOp__strm1_data_valid =  sti__stOp__lane12_strm1_data_valid    ;
  // Lane 13, Stream 1
  assign stOp__sti__lane13_strm1_ready             =  stOp_lane[13].stOp__sti__strm1_ready  ;
  assign stOp_lane[13].sti__stOp__strm1_cntl       =  sti__stOp__lane13_strm1_cntl          ;
  assign stOp_lane[13].sti__stOp__strm1_data       =  sti__stOp__lane13_strm1_data          ;
  assign stOp_lane[13].sti__stOp__strm1_data_valid =  sti__stOp__lane13_strm1_data_valid    ;
  // Lane 14, Stream 1
  assign stOp__sti__lane14_strm1_ready             =  stOp_lane[14].stOp__sti__strm1_ready  ;
  assign stOp_lane[14].sti__stOp__strm1_cntl       =  sti__stOp__lane14_strm1_cntl          ;
  assign stOp_lane[14].sti__stOp__strm1_data       =  sti__stOp__lane14_strm1_data          ;
  assign stOp_lane[14].sti__stOp__strm1_data_valid =  sti__stOp__lane14_strm1_data_valid    ;
  // Lane 15, Stream 1
  assign stOp__sti__lane15_strm1_ready             =  stOp_lane[15].stOp__sti__strm1_ready  ;
  assign stOp_lane[15].sti__stOp__strm1_cntl       =  sti__stOp__lane15_strm1_cntl          ;
  assign stOp_lane[15].sti__stOp__strm1_data       =  sti__stOp__lane15_strm1_data          ;
  assign stOp_lane[15].sti__stOp__strm1_data_valid =  sti__stOp__lane15_strm1_data_valid    ;
  // Lane 16, Stream 1
  assign stOp__sti__lane16_strm1_ready             =  stOp_lane[16].stOp__sti__strm1_ready  ;
  assign stOp_lane[16].sti__stOp__strm1_cntl       =  sti__stOp__lane16_strm1_cntl          ;
  assign stOp_lane[16].sti__stOp__strm1_data       =  sti__stOp__lane16_strm1_data          ;
  assign stOp_lane[16].sti__stOp__strm1_data_valid =  sti__stOp__lane16_strm1_data_valid    ;
  // Lane 17, Stream 1
  assign stOp__sti__lane17_strm1_ready             =  stOp_lane[17].stOp__sti__strm1_ready  ;
  assign stOp_lane[17].sti__stOp__strm1_cntl       =  sti__stOp__lane17_strm1_cntl          ;
  assign stOp_lane[17].sti__stOp__strm1_data       =  sti__stOp__lane17_strm1_data          ;
  assign stOp_lane[17].sti__stOp__strm1_data_valid =  sti__stOp__lane17_strm1_data_valid    ;
  // Lane 18, Stream 1
  assign stOp__sti__lane18_strm1_ready             =  stOp_lane[18].stOp__sti__strm1_ready  ;
  assign stOp_lane[18].sti__stOp__strm1_cntl       =  sti__stOp__lane18_strm1_cntl          ;
  assign stOp_lane[18].sti__stOp__strm1_data       =  sti__stOp__lane18_strm1_data          ;
  assign stOp_lane[18].sti__stOp__strm1_data_valid =  sti__stOp__lane18_strm1_data_valid    ;
  // Lane 19, Stream 1
  assign stOp__sti__lane19_strm1_ready             =  stOp_lane[19].stOp__sti__strm1_ready  ;
  assign stOp_lane[19].sti__stOp__strm1_cntl       =  sti__stOp__lane19_strm1_cntl          ;
  assign stOp_lane[19].sti__stOp__strm1_data       =  sti__stOp__lane19_strm1_data          ;
  assign stOp_lane[19].sti__stOp__strm1_data_valid =  sti__stOp__lane19_strm1_data_valid    ;
  // Lane 20, Stream 1
  assign stOp__sti__lane20_strm1_ready             =  stOp_lane[20].stOp__sti__strm1_ready  ;
  assign stOp_lane[20].sti__stOp__strm1_cntl       =  sti__stOp__lane20_strm1_cntl          ;
  assign stOp_lane[20].sti__stOp__strm1_data       =  sti__stOp__lane20_strm1_data          ;
  assign stOp_lane[20].sti__stOp__strm1_data_valid =  sti__stOp__lane20_strm1_data_valid    ;
  // Lane 21, Stream 1
  assign stOp__sti__lane21_strm1_ready             =  stOp_lane[21].stOp__sti__strm1_ready  ;
  assign stOp_lane[21].sti__stOp__strm1_cntl       =  sti__stOp__lane21_strm1_cntl          ;
  assign stOp_lane[21].sti__stOp__strm1_data       =  sti__stOp__lane21_strm1_data          ;
  assign stOp_lane[21].sti__stOp__strm1_data_valid =  sti__stOp__lane21_strm1_data_valid    ;
  // Lane 22, Stream 1
  assign stOp__sti__lane22_strm1_ready             =  stOp_lane[22].stOp__sti__strm1_ready  ;
  assign stOp_lane[22].sti__stOp__strm1_cntl       =  sti__stOp__lane22_strm1_cntl          ;
  assign stOp_lane[22].sti__stOp__strm1_data       =  sti__stOp__lane22_strm1_data          ;
  assign stOp_lane[22].sti__stOp__strm1_data_valid =  sti__stOp__lane22_strm1_data_valid    ;
  // Lane 23, Stream 1
  assign stOp__sti__lane23_strm1_ready             =  stOp_lane[23].stOp__sti__strm1_ready  ;
  assign stOp_lane[23].sti__stOp__strm1_cntl       =  sti__stOp__lane23_strm1_cntl          ;
  assign stOp_lane[23].sti__stOp__strm1_data       =  sti__stOp__lane23_strm1_data          ;
  assign stOp_lane[23].sti__stOp__strm1_data_valid =  sti__stOp__lane23_strm1_data_valid    ;
  // Lane 24, Stream 1
  assign stOp__sti__lane24_strm1_ready             =  stOp_lane[24].stOp__sti__strm1_ready  ;
  assign stOp_lane[24].sti__stOp__strm1_cntl       =  sti__stOp__lane24_strm1_cntl          ;
  assign stOp_lane[24].sti__stOp__strm1_data       =  sti__stOp__lane24_strm1_data          ;
  assign stOp_lane[24].sti__stOp__strm1_data_valid =  sti__stOp__lane24_strm1_data_valid    ;
  // Lane 25, Stream 1
  assign stOp__sti__lane25_strm1_ready             =  stOp_lane[25].stOp__sti__strm1_ready  ;
  assign stOp_lane[25].sti__stOp__strm1_cntl       =  sti__stOp__lane25_strm1_cntl          ;
  assign stOp_lane[25].sti__stOp__strm1_data       =  sti__stOp__lane25_strm1_data          ;
  assign stOp_lane[25].sti__stOp__strm1_data_valid =  sti__stOp__lane25_strm1_data_valid    ;
  // Lane 26, Stream 1
  assign stOp__sti__lane26_strm1_ready             =  stOp_lane[26].stOp__sti__strm1_ready  ;
  assign stOp_lane[26].sti__stOp__strm1_cntl       =  sti__stOp__lane26_strm1_cntl          ;
  assign stOp_lane[26].sti__stOp__strm1_data       =  sti__stOp__lane26_strm1_data          ;
  assign stOp_lane[26].sti__stOp__strm1_data_valid =  sti__stOp__lane26_strm1_data_valid    ;
  // Lane 27, Stream 1
  assign stOp__sti__lane27_strm1_ready             =  stOp_lane[27].stOp__sti__strm1_ready  ;
  assign stOp_lane[27].sti__stOp__strm1_cntl       =  sti__stOp__lane27_strm1_cntl          ;
  assign stOp_lane[27].sti__stOp__strm1_data       =  sti__stOp__lane27_strm1_data          ;
  assign stOp_lane[27].sti__stOp__strm1_data_valid =  sti__stOp__lane27_strm1_data_valid    ;
  // Lane 28, Stream 1
  assign stOp__sti__lane28_strm1_ready             =  stOp_lane[28].stOp__sti__strm1_ready  ;
  assign stOp_lane[28].sti__stOp__strm1_cntl       =  sti__stOp__lane28_strm1_cntl          ;
  assign stOp_lane[28].sti__stOp__strm1_data       =  sti__stOp__lane28_strm1_data          ;
  assign stOp_lane[28].sti__stOp__strm1_data_valid =  sti__stOp__lane28_strm1_data_valid    ;
  // Lane 29, Stream 1
  assign stOp__sti__lane29_strm1_ready             =  stOp_lane[29].stOp__sti__strm1_ready  ;
  assign stOp_lane[29].sti__stOp__strm1_cntl       =  sti__stOp__lane29_strm1_cntl          ;
  assign stOp_lane[29].sti__stOp__strm1_data       =  sti__stOp__lane29_strm1_data          ;
  assign stOp_lane[29].sti__stOp__strm1_data_valid =  sti__stOp__lane29_strm1_data_valid    ;
  // Lane 30, Stream 1
  assign stOp__sti__lane30_strm1_ready             =  stOp_lane[30].stOp__sti__strm1_ready  ;
  assign stOp_lane[30].sti__stOp__strm1_cntl       =  sti__stOp__lane30_strm1_cntl          ;
  assign stOp_lane[30].sti__stOp__strm1_data       =  sti__stOp__lane30_strm1_data          ;
  assign stOp_lane[30].sti__stOp__strm1_data_valid =  sti__stOp__lane30_strm1_data_valid    ;
  // Lane 31, Stream 1
  assign stOp__sti__lane31_strm1_ready             =  stOp_lane[31].stOp__sti__strm1_ready  ;
  assign stOp_lane[31].sti__stOp__strm1_cntl       =  sti__stOp__lane31_strm1_cntl          ;
  assign stOp_lane[31].sti__stOp__strm1_data       =  sti__stOp__lane31_strm1_data          ;
  assign stOp_lane[31].sti__stOp__strm1_data_valid =  sti__stOp__lane31_strm1_data_valid    ;
