
//------------------------------------------------
// MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_LOCAL_INPUT_QUEUE_CONTROL_STATE width
//------------------------------------------------
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_STATE_MSB            16
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_STATE_LSB            0
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_STATE_SIZE           (`MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_STATE_MSB - `MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_STATE_LSB +1)
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_STATE_RANGE           `MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_STATE_MSB : `MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_STATE_LSB

//------------------------------------------------------------------------------------------------
//------------------------------------------------
// MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL state machine states
//------------------------------------------------

`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_WAIT        17'd1
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_WAIT_START_LOCAL  17'd2
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_TRANSFER_LOCAL  17'd4
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_ACK_LOCAL   17'd8
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_WAIT_START_PORT0  17'd16
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_TRANSFER_PORT0  17'd32
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_ACK_PORT0   17'd64
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_WAIT_START_PORT1  17'd128
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_TRANSFER_PORT1  17'd256
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_ACK_PORT1   17'd512
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_WAIT_START_PORT2  17'd1024
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_TRANSFER_PORT2  17'd2048
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_ACK_PORT2   17'd4096
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_WAIT_START_PORT3  17'd8192
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_TRANSFER_PORT3  17'd16384
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_ACK_PORT3   17'd32768
`define MGR_NOC_CONT_NOC_PORT_OUTPUT_CNTL_ERR   17'd65536