

            // ##################################################
            // DMA Stream Destination addresses

            // Stream 0 Destination address
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [0] = 32'b000000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [1] = 32'b000000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [2] = 32'b000000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [3] = 32'b000000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [4] = 32'b000000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [5] = 32'b000000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [6] = 32'b000000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [7] = 32'b000000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [8] = 32'b000000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [9] = 32'b000000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [10] = 32'b000000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [11] = 32'b000000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [12] = 32'b000000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [13] = 32'b000000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [14] = 32'b000000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [15] = 32'b000000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [16] = 32'b000000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [17] = 32'b000000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [18] = 32'b000000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [19] = 32'b000000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [20] = 32'b000000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [21] = 32'b000000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [22] = 32'b000000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [23] = 32'b000000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [24] = 32'b000000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [25] = 32'b000000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [26] = 32'b000000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [27] = 32'b000000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [28] = 32'b000000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [29] = 32'b000000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [30] = 32'b000000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [31] = 32'b000000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [0] = 32'b000000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [1] = 32'b000000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [2] = 32'b000000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [3] = 32'b000000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [4] = 32'b000000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [5] = 32'b000000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [6] = 32'b000000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [7] = 32'b000000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [8] = 32'b000000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [9] = 32'b000000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [10] = 32'b000000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [11] = 32'b000000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [12] = 32'b000000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [13] = 32'b000000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [14] = 32'b000000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [15] = 32'b000000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [16] = 32'b000000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [17] = 32'b000000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [18] = 32'b000000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [19] = 32'b000000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [20] = 32'b000000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [21] = 32'b000000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [22] = 32'b000000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [23] = 32'b000000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [24] = 32'b000000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [25] = 32'b000000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [26] = 32'b000000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [27] = 32'b000000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [28] = 32'b000000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [29] = 32'b000000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [30] = 32'b000000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [31] = 32'b000000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [0] = 32'b000001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [1] = 32'b000001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [2] = 32'b000001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [3] = 32'b000001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [4] = 32'b000001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [5] = 32'b000001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [6] = 32'b000001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [7] = 32'b000001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [8] = 32'b000001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [9] = 32'b000001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [10] = 32'b000001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [11] = 32'b000001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [12] = 32'b000001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [13] = 32'b000001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [14] = 32'b000001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [15] = 32'b000001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [16] = 32'b000001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [17] = 32'b000001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [18] = 32'b000001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [19] = 32'b000001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [20] = 32'b000001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [21] = 32'b000001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [22] = 32'b000001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [23] = 32'b000001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [24] = 32'b000001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [25] = 32'b000001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [26] = 32'b000001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [27] = 32'b000001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [28] = 32'b000001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [29] = 32'b000001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [30] = 32'b000001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [31] = 32'b000001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [0] = 32'b000001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [1] = 32'b000001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [2] = 32'b000001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [3] = 32'b000001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [4] = 32'b000001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [5] = 32'b000001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [6] = 32'b000001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [7] = 32'b000001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [8] = 32'b000001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [9] = 32'b000001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [10] = 32'b000001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [11] = 32'b000001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [12] = 32'b000001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [13] = 32'b000001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [14] = 32'b000001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [15] = 32'b000001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [16] = 32'b000001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [17] = 32'b000001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [18] = 32'b000001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [19] = 32'b000001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [20] = 32'b000001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [21] = 32'b000001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [22] = 32'b000001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [23] = 32'b000001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [24] = 32'b000001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [25] = 32'b000001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [26] = 32'b000001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [27] = 32'b000001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [28] = 32'b000001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [29] = 32'b000001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [30] = 32'b000001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [31] = 32'b000001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [0] = 32'b000010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [1] = 32'b000010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [2] = 32'b000010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [3] = 32'b000010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [4] = 32'b000010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [5] = 32'b000010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [6] = 32'b000010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [7] = 32'b000010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [8] = 32'b000010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [9] = 32'b000010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [10] = 32'b000010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [11] = 32'b000010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [12] = 32'b000010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [13] = 32'b000010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [14] = 32'b000010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [15] = 32'b000010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [16] = 32'b000010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [17] = 32'b000010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [18] = 32'b000010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [19] = 32'b000010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [20] = 32'b000010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [21] = 32'b000010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [22] = 32'b000010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [23] = 32'b000010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [24] = 32'b000010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [25] = 32'b000010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [26] = 32'b000010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [27] = 32'b000010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [28] = 32'b000010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [29] = 32'b000010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [30] = 32'b000010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [31] = 32'b000010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [0] = 32'b000010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [1] = 32'b000010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [2] = 32'b000010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [3] = 32'b000010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [4] = 32'b000010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [5] = 32'b000010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [6] = 32'b000010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [7] = 32'b000010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [8] = 32'b000010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [9] = 32'b000010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [10] = 32'b000010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [11] = 32'b000010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [12] = 32'b000010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [13] = 32'b000010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [14] = 32'b000010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [15] = 32'b000010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [16] = 32'b000010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [17] = 32'b000010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [18] = 32'b000010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [19] = 32'b000010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [20] = 32'b000010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [21] = 32'b000010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [22] = 32'b000010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [23] = 32'b000010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [24] = 32'b000010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [25] = 32'b000010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [26] = 32'b000010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [27] = 32'b000010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [28] = 32'b000010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [29] = 32'b000010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [30] = 32'b000010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [31] = 32'b000010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [0] = 32'b000011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [1] = 32'b000011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [2] = 32'b000011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [3] = 32'b000011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [4] = 32'b000011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [5] = 32'b000011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [6] = 32'b000011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [7] = 32'b000011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [8] = 32'b000011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [9] = 32'b000011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [10] = 32'b000011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [11] = 32'b000011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [12] = 32'b000011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [13] = 32'b000011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [14] = 32'b000011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [15] = 32'b000011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [16] = 32'b000011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [17] = 32'b000011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [18] = 32'b000011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [19] = 32'b000011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [20] = 32'b000011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [21] = 32'b000011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [22] = 32'b000011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [23] = 32'b000011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [24] = 32'b000011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [25] = 32'b000011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [26] = 32'b000011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [27] = 32'b000011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [28] = 32'b000011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [29] = 32'b000011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [30] = 32'b000011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [31] = 32'b000011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [0] = 32'b000011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [1] = 32'b000011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [2] = 32'b000011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [3] = 32'b000011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [4] = 32'b000011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [5] = 32'b000011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [6] = 32'b000011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [7] = 32'b000011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [8] = 32'b000011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [9] = 32'b000011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [10] = 32'b000011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [11] = 32'b000011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [12] = 32'b000011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [13] = 32'b000011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [14] = 32'b000011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [15] = 32'b000011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [16] = 32'b000011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [17] = 32'b000011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [18] = 32'b000011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [19] = 32'b000011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [20] = 32'b000011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [21] = 32'b000011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [22] = 32'b000011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [23] = 32'b000011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [24] = 32'b000011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [25] = 32'b000011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [26] = 32'b000011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [27] = 32'b000011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [28] = 32'b000011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [29] = 32'b000011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [30] = 32'b000011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [31] = 32'b000011_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [0] = 32'b000100_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [1] = 32'b000100_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [2] = 32'b000100_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [3] = 32'b000100_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [4] = 32'b000100_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [5] = 32'b000100_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [6] = 32'b000100_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [7] = 32'b000100_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [8] = 32'b000100_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [9] = 32'b000100_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [10] = 32'b000100_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [11] = 32'b000100_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [12] = 32'b000100_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [13] = 32'b000100_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [14] = 32'b000100_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [15] = 32'b000100_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [16] = 32'b000100_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [17] = 32'b000100_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [18] = 32'b000100_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [19] = 32'b000100_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [20] = 32'b000100_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [21] = 32'b000100_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [22] = 32'b000100_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [23] = 32'b000100_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [24] = 32'b000100_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [25] = 32'b000100_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [26] = 32'b000100_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [27] = 32'b000100_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [28] = 32'b000100_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [29] = 32'b000100_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [30] = 32'b000100_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r134 [31] = 32'b000100_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [0] = 32'b000100_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [1] = 32'b000100_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [2] = 32'b000100_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [3] = 32'b000100_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [4] = 32'b000100_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [5] = 32'b000100_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [6] = 32'b000100_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [7] = 32'b000100_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [8] = 32'b000100_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [9] = 32'b000100_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [10] = 32'b000100_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [11] = 32'b000100_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [12] = 32'b000100_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [13] = 32'b000100_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [14] = 32'b000100_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [15] = 32'b000100_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [16] = 32'b000100_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [17] = 32'b000100_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [18] = 32'b000100_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [19] = 32'b000100_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [20] = 32'b000100_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [21] = 32'b000100_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [22] = 32'b000100_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [23] = 32'b000100_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [24] = 32'b000100_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [25] = 32'b000100_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [26] = 32'b000100_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [27] = 32'b000100_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [28] = 32'b000100_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [29] = 32'b000100_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [30] = 32'b000100_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r135 [31] = 32'b000100_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [0] = 32'b000101_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [1] = 32'b000101_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [2] = 32'b000101_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [3] = 32'b000101_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [4] = 32'b000101_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [5] = 32'b000101_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [6] = 32'b000101_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [7] = 32'b000101_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [8] = 32'b000101_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [9] = 32'b000101_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [10] = 32'b000101_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [11] = 32'b000101_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [12] = 32'b000101_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [13] = 32'b000101_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [14] = 32'b000101_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [15] = 32'b000101_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [16] = 32'b000101_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [17] = 32'b000101_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [18] = 32'b000101_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [19] = 32'b000101_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [20] = 32'b000101_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [21] = 32'b000101_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [22] = 32'b000101_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [23] = 32'b000101_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [24] = 32'b000101_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [25] = 32'b000101_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [26] = 32'b000101_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [27] = 32'b000101_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [28] = 32'b000101_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [29] = 32'b000101_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [30] = 32'b000101_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r134 [31] = 32'b000101_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [0] = 32'b000101_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [1] = 32'b000101_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [2] = 32'b000101_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [3] = 32'b000101_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [4] = 32'b000101_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [5] = 32'b000101_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [6] = 32'b000101_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [7] = 32'b000101_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [8] = 32'b000101_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [9] = 32'b000101_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [10] = 32'b000101_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [11] = 32'b000101_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [12] = 32'b000101_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [13] = 32'b000101_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [14] = 32'b000101_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [15] = 32'b000101_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [16] = 32'b000101_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [17] = 32'b000101_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [18] = 32'b000101_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [19] = 32'b000101_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [20] = 32'b000101_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [21] = 32'b000101_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [22] = 32'b000101_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [23] = 32'b000101_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [24] = 32'b000101_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [25] = 32'b000101_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [26] = 32'b000101_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [27] = 32'b000101_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [28] = 32'b000101_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [29] = 32'b000101_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [30] = 32'b000101_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r135 [31] = 32'b000101_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [0] = 32'b000110_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [1] = 32'b000110_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [2] = 32'b000110_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [3] = 32'b000110_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [4] = 32'b000110_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [5] = 32'b000110_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [6] = 32'b000110_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [7] = 32'b000110_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [8] = 32'b000110_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [9] = 32'b000110_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [10] = 32'b000110_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [11] = 32'b000110_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [12] = 32'b000110_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [13] = 32'b000110_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [14] = 32'b000110_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [15] = 32'b000110_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [16] = 32'b000110_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [17] = 32'b000110_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [18] = 32'b000110_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [19] = 32'b000110_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [20] = 32'b000110_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [21] = 32'b000110_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [22] = 32'b000110_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [23] = 32'b000110_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [24] = 32'b000110_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [25] = 32'b000110_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [26] = 32'b000110_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [27] = 32'b000110_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [28] = 32'b000110_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [29] = 32'b000110_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [30] = 32'b000110_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r134 [31] = 32'b000110_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [0] = 32'b000110_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [1] = 32'b000110_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [2] = 32'b000110_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [3] = 32'b000110_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [4] = 32'b000110_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [5] = 32'b000110_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [6] = 32'b000110_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [7] = 32'b000110_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [8] = 32'b000110_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [9] = 32'b000110_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [10] = 32'b000110_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [11] = 32'b000110_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [12] = 32'b000110_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [13] = 32'b000110_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [14] = 32'b000110_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [15] = 32'b000110_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [16] = 32'b000110_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [17] = 32'b000110_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [18] = 32'b000110_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [19] = 32'b000110_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [20] = 32'b000110_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [21] = 32'b000110_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [22] = 32'b000110_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [23] = 32'b000110_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [24] = 32'b000110_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [25] = 32'b000110_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [26] = 32'b000110_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [27] = 32'b000110_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [28] = 32'b000110_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [29] = 32'b000110_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [30] = 32'b000110_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r135 [31] = 32'b000110_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [0] = 32'b000111_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [1] = 32'b000111_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [2] = 32'b000111_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [3] = 32'b000111_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [4] = 32'b000111_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [5] = 32'b000111_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [6] = 32'b000111_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [7] = 32'b000111_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [8] = 32'b000111_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [9] = 32'b000111_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [10] = 32'b000111_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [11] = 32'b000111_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [12] = 32'b000111_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [13] = 32'b000111_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [14] = 32'b000111_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [15] = 32'b000111_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [16] = 32'b000111_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [17] = 32'b000111_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [18] = 32'b000111_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [19] = 32'b000111_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [20] = 32'b000111_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [21] = 32'b000111_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [22] = 32'b000111_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [23] = 32'b000111_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [24] = 32'b000111_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [25] = 32'b000111_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [26] = 32'b000111_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [27] = 32'b000111_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [28] = 32'b000111_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [29] = 32'b000111_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [30] = 32'b000111_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r134 [31] = 32'b000111_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [0] = 32'b000111_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [1] = 32'b000111_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [2] = 32'b000111_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [3] = 32'b000111_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [4] = 32'b000111_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [5] = 32'b000111_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [6] = 32'b000111_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [7] = 32'b000111_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [8] = 32'b000111_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [9] = 32'b000111_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [10] = 32'b000111_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [11] = 32'b000111_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [12] = 32'b000111_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [13] = 32'b000111_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [14] = 32'b000111_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [15] = 32'b000111_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [16] = 32'b000111_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [17] = 32'b000111_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [18] = 32'b000111_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [19] = 32'b000111_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [20] = 32'b000111_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [21] = 32'b000111_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [22] = 32'b000111_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [23] = 32'b000111_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [24] = 32'b000111_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [25] = 32'b000111_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [26] = 32'b000111_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [27] = 32'b000111_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [28] = 32'b000111_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [29] = 32'b000111_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [30] = 32'b000111_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r135 [31] = 32'b000111_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [0] = 32'b001000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [1] = 32'b001000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [2] = 32'b001000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [3] = 32'b001000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [4] = 32'b001000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [5] = 32'b001000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [6] = 32'b001000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [7] = 32'b001000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [8] = 32'b001000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [9] = 32'b001000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [10] = 32'b001000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [11] = 32'b001000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [12] = 32'b001000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [13] = 32'b001000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [14] = 32'b001000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [15] = 32'b001000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [16] = 32'b001000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [17] = 32'b001000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [18] = 32'b001000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [19] = 32'b001000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [20] = 32'b001000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [21] = 32'b001000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [22] = 32'b001000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [23] = 32'b001000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [24] = 32'b001000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [25] = 32'b001000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [26] = 32'b001000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [27] = 32'b001000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [28] = 32'b001000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [29] = 32'b001000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [30] = 32'b001000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r134 [31] = 32'b001000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [0] = 32'b001000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [1] = 32'b001000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [2] = 32'b001000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [3] = 32'b001000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [4] = 32'b001000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [5] = 32'b001000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [6] = 32'b001000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [7] = 32'b001000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [8] = 32'b001000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [9] = 32'b001000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [10] = 32'b001000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [11] = 32'b001000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [12] = 32'b001000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [13] = 32'b001000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [14] = 32'b001000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [15] = 32'b001000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [16] = 32'b001000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [17] = 32'b001000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [18] = 32'b001000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [19] = 32'b001000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [20] = 32'b001000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [21] = 32'b001000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [22] = 32'b001000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [23] = 32'b001000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [24] = 32'b001000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [25] = 32'b001000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [26] = 32'b001000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [27] = 32'b001000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [28] = 32'b001000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [29] = 32'b001000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [30] = 32'b001000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r135 [31] = 32'b001000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [0] = 32'b001001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [1] = 32'b001001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [2] = 32'b001001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [3] = 32'b001001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [4] = 32'b001001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [5] = 32'b001001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [6] = 32'b001001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [7] = 32'b001001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [8] = 32'b001001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [9] = 32'b001001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [10] = 32'b001001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [11] = 32'b001001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [12] = 32'b001001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [13] = 32'b001001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [14] = 32'b001001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [15] = 32'b001001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [16] = 32'b001001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [17] = 32'b001001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [18] = 32'b001001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [19] = 32'b001001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [20] = 32'b001001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [21] = 32'b001001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [22] = 32'b001001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [23] = 32'b001001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [24] = 32'b001001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [25] = 32'b001001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [26] = 32'b001001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [27] = 32'b001001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [28] = 32'b001001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [29] = 32'b001001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [30] = 32'b001001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r134 [31] = 32'b001001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [0] = 32'b001001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [1] = 32'b001001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [2] = 32'b001001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [3] = 32'b001001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [4] = 32'b001001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [5] = 32'b001001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [6] = 32'b001001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [7] = 32'b001001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [8] = 32'b001001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [9] = 32'b001001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [10] = 32'b001001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [11] = 32'b001001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [12] = 32'b001001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [13] = 32'b001001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [14] = 32'b001001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [15] = 32'b001001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [16] = 32'b001001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [17] = 32'b001001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [18] = 32'b001001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [19] = 32'b001001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [20] = 32'b001001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [21] = 32'b001001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [22] = 32'b001001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [23] = 32'b001001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [24] = 32'b001001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [25] = 32'b001001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [26] = 32'b001001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [27] = 32'b001001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [28] = 32'b001001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [29] = 32'b001001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [30] = 32'b001001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r135 [31] = 32'b001001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [0] = 32'b001010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [1] = 32'b001010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [2] = 32'b001010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [3] = 32'b001010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [4] = 32'b001010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [5] = 32'b001010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [6] = 32'b001010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [7] = 32'b001010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [8] = 32'b001010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [9] = 32'b001010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [10] = 32'b001010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [11] = 32'b001010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [12] = 32'b001010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [13] = 32'b001010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [14] = 32'b001010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [15] = 32'b001010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [16] = 32'b001010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [17] = 32'b001010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [18] = 32'b001010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [19] = 32'b001010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [20] = 32'b001010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [21] = 32'b001010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [22] = 32'b001010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [23] = 32'b001010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [24] = 32'b001010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [25] = 32'b001010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [26] = 32'b001010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [27] = 32'b001010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [28] = 32'b001010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [29] = 32'b001010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [30] = 32'b001010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r134 [31] = 32'b001010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [0] = 32'b001010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [1] = 32'b001010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [2] = 32'b001010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [3] = 32'b001010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [4] = 32'b001010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [5] = 32'b001010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [6] = 32'b001010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [7] = 32'b001010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [8] = 32'b001010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [9] = 32'b001010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [10] = 32'b001010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [11] = 32'b001010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [12] = 32'b001010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [13] = 32'b001010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [14] = 32'b001010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [15] = 32'b001010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [16] = 32'b001010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [17] = 32'b001010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [18] = 32'b001010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [19] = 32'b001010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [20] = 32'b001010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [21] = 32'b001010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [22] = 32'b001010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [23] = 32'b001010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [24] = 32'b001010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [25] = 32'b001010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [26] = 32'b001010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [27] = 32'b001010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [28] = 32'b001010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [29] = 32'b001010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [30] = 32'b001010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r135 [31] = 32'b001010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [0] = 32'b001011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [1] = 32'b001011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [2] = 32'b001011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [3] = 32'b001011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [4] = 32'b001011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [5] = 32'b001011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [6] = 32'b001011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [7] = 32'b001011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [8] = 32'b001011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [9] = 32'b001011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [10] = 32'b001011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [11] = 32'b001011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [12] = 32'b001011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [13] = 32'b001011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [14] = 32'b001011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [15] = 32'b001011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [16] = 32'b001011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [17] = 32'b001011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [18] = 32'b001011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [19] = 32'b001011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [20] = 32'b001011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [21] = 32'b001011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [22] = 32'b001011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [23] = 32'b001011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [24] = 32'b001011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [25] = 32'b001011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [26] = 32'b001011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [27] = 32'b001011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [28] = 32'b001011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [29] = 32'b001011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [30] = 32'b001011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r134 [31] = 32'b001011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [0] = 32'b001011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [1] = 32'b001011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [2] = 32'b001011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [3] = 32'b001011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [4] = 32'b001011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [5] = 32'b001011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [6] = 32'b001011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [7] = 32'b001011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [8] = 32'b001011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [9] = 32'b001011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [10] = 32'b001011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [11] = 32'b001011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [12] = 32'b001011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [13] = 32'b001011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [14] = 32'b001011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [15] = 32'b001011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [16] = 32'b001011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [17] = 32'b001011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [18] = 32'b001011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [19] = 32'b001011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [20] = 32'b001011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [21] = 32'b001011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [22] = 32'b001011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [23] = 32'b001011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [24] = 32'b001011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [25] = 32'b001011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [26] = 32'b001011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [27] = 32'b001011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [28] = 32'b001011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [29] = 32'b001011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [30] = 32'b001011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r135 [31] = 32'b001011_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [0] = 32'b001100_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [1] = 32'b001100_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [2] = 32'b001100_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [3] = 32'b001100_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [4] = 32'b001100_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [5] = 32'b001100_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [6] = 32'b001100_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [7] = 32'b001100_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [8] = 32'b001100_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [9] = 32'b001100_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [10] = 32'b001100_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [11] = 32'b001100_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [12] = 32'b001100_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [13] = 32'b001100_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [14] = 32'b001100_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [15] = 32'b001100_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [16] = 32'b001100_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [17] = 32'b001100_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [18] = 32'b001100_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [19] = 32'b001100_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [20] = 32'b001100_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [21] = 32'b001100_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [22] = 32'b001100_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [23] = 32'b001100_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [24] = 32'b001100_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [25] = 32'b001100_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [26] = 32'b001100_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [27] = 32'b001100_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [28] = 32'b001100_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [29] = 32'b001100_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [30] = 32'b001100_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r134 [31] = 32'b001100_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [0] = 32'b001100_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [1] = 32'b001100_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [2] = 32'b001100_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [3] = 32'b001100_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [4] = 32'b001100_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [5] = 32'b001100_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [6] = 32'b001100_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [7] = 32'b001100_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [8] = 32'b001100_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [9] = 32'b001100_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [10] = 32'b001100_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [11] = 32'b001100_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [12] = 32'b001100_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [13] = 32'b001100_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [14] = 32'b001100_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [15] = 32'b001100_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [16] = 32'b001100_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [17] = 32'b001100_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [18] = 32'b001100_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [19] = 32'b001100_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [20] = 32'b001100_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [21] = 32'b001100_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [22] = 32'b001100_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [23] = 32'b001100_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [24] = 32'b001100_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [25] = 32'b001100_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [26] = 32'b001100_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [27] = 32'b001100_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [28] = 32'b001100_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [29] = 32'b001100_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [30] = 32'b001100_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r135 [31] = 32'b001100_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [0] = 32'b001101_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [1] = 32'b001101_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [2] = 32'b001101_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [3] = 32'b001101_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [4] = 32'b001101_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [5] = 32'b001101_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [6] = 32'b001101_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [7] = 32'b001101_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [8] = 32'b001101_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [9] = 32'b001101_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [10] = 32'b001101_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [11] = 32'b001101_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [12] = 32'b001101_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [13] = 32'b001101_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [14] = 32'b001101_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [15] = 32'b001101_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [16] = 32'b001101_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [17] = 32'b001101_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [18] = 32'b001101_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [19] = 32'b001101_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [20] = 32'b001101_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [21] = 32'b001101_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [22] = 32'b001101_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [23] = 32'b001101_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [24] = 32'b001101_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [25] = 32'b001101_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [26] = 32'b001101_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [27] = 32'b001101_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [28] = 32'b001101_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [29] = 32'b001101_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [30] = 32'b001101_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r134 [31] = 32'b001101_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [0] = 32'b001101_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [1] = 32'b001101_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [2] = 32'b001101_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [3] = 32'b001101_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [4] = 32'b001101_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [5] = 32'b001101_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [6] = 32'b001101_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [7] = 32'b001101_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [8] = 32'b001101_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [9] = 32'b001101_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [10] = 32'b001101_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [11] = 32'b001101_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [12] = 32'b001101_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [13] = 32'b001101_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [14] = 32'b001101_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [15] = 32'b001101_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [16] = 32'b001101_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [17] = 32'b001101_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [18] = 32'b001101_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [19] = 32'b001101_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [20] = 32'b001101_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [21] = 32'b001101_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [22] = 32'b001101_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [23] = 32'b001101_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [24] = 32'b001101_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [25] = 32'b001101_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [26] = 32'b001101_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [27] = 32'b001101_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [28] = 32'b001101_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [29] = 32'b001101_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [30] = 32'b001101_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r135 [31] = 32'b001101_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [0] = 32'b001110_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [1] = 32'b001110_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [2] = 32'b001110_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [3] = 32'b001110_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [4] = 32'b001110_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [5] = 32'b001110_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [6] = 32'b001110_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [7] = 32'b001110_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [8] = 32'b001110_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [9] = 32'b001110_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [10] = 32'b001110_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [11] = 32'b001110_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [12] = 32'b001110_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [13] = 32'b001110_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [14] = 32'b001110_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [15] = 32'b001110_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [16] = 32'b001110_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [17] = 32'b001110_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [18] = 32'b001110_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [19] = 32'b001110_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [20] = 32'b001110_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [21] = 32'b001110_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [22] = 32'b001110_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [23] = 32'b001110_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [24] = 32'b001110_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [25] = 32'b001110_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [26] = 32'b001110_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [27] = 32'b001110_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [28] = 32'b001110_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [29] = 32'b001110_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [30] = 32'b001110_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r134 [31] = 32'b001110_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [0] = 32'b001110_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [1] = 32'b001110_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [2] = 32'b001110_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [3] = 32'b001110_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [4] = 32'b001110_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [5] = 32'b001110_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [6] = 32'b001110_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [7] = 32'b001110_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [8] = 32'b001110_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [9] = 32'b001110_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [10] = 32'b001110_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [11] = 32'b001110_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [12] = 32'b001110_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [13] = 32'b001110_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [14] = 32'b001110_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [15] = 32'b001110_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [16] = 32'b001110_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [17] = 32'b001110_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [18] = 32'b001110_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [19] = 32'b001110_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [20] = 32'b001110_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [21] = 32'b001110_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [22] = 32'b001110_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [23] = 32'b001110_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [24] = 32'b001110_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [25] = 32'b001110_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [26] = 32'b001110_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [27] = 32'b001110_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [28] = 32'b001110_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [29] = 32'b001110_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [30] = 32'b001110_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r135 [31] = 32'b001110_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [0] = 32'b001111_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [1] = 32'b001111_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [2] = 32'b001111_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [3] = 32'b001111_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [4] = 32'b001111_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [5] = 32'b001111_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [6] = 32'b001111_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [7] = 32'b001111_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [8] = 32'b001111_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [9] = 32'b001111_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [10] = 32'b001111_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [11] = 32'b001111_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [12] = 32'b001111_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [13] = 32'b001111_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [14] = 32'b001111_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [15] = 32'b001111_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [16] = 32'b001111_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [17] = 32'b001111_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [18] = 32'b001111_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [19] = 32'b001111_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [20] = 32'b001111_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [21] = 32'b001111_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [22] = 32'b001111_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [23] = 32'b001111_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [24] = 32'b001111_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [25] = 32'b001111_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [26] = 32'b001111_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [27] = 32'b001111_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [28] = 32'b001111_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [29] = 32'b001111_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [30] = 32'b001111_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r134 [31] = 32'b001111_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [0] = 32'b001111_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [1] = 32'b001111_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [2] = 32'b001111_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [3] = 32'b001111_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [4] = 32'b001111_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [5] = 32'b001111_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [6] = 32'b001111_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [7] = 32'b001111_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [8] = 32'b001111_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [9] = 32'b001111_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [10] = 32'b001111_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [11] = 32'b001111_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [12] = 32'b001111_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [13] = 32'b001111_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [14] = 32'b001111_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [15] = 32'b001111_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [16] = 32'b001111_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [17] = 32'b001111_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [18] = 32'b001111_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [19] = 32'b001111_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [20] = 32'b001111_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [21] = 32'b001111_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [22] = 32'b001111_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [23] = 32'b001111_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [24] = 32'b001111_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [25] = 32'b001111_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [26] = 32'b001111_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [27] = 32'b001111_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [28] = 32'b001111_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [29] = 32'b001111_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [30] = 32'b001111_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r135 [31] = 32'b001111_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [0] = 32'b010000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [1] = 32'b010000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [2] = 32'b010000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [3] = 32'b010000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [4] = 32'b010000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [5] = 32'b010000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [6] = 32'b010000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [7] = 32'b010000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [8] = 32'b010000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [9] = 32'b010000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [10] = 32'b010000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [11] = 32'b010000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [12] = 32'b010000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [13] = 32'b010000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [14] = 32'b010000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [15] = 32'b010000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [16] = 32'b010000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [17] = 32'b010000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [18] = 32'b010000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [19] = 32'b010000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [20] = 32'b010000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [21] = 32'b010000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [22] = 32'b010000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [23] = 32'b010000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [24] = 32'b010000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [25] = 32'b010000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [26] = 32'b010000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [27] = 32'b010000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [28] = 32'b010000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [29] = 32'b010000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [30] = 32'b010000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r134 [31] = 32'b010000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [0] = 32'b010000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [1] = 32'b010000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [2] = 32'b010000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [3] = 32'b010000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [4] = 32'b010000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [5] = 32'b010000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [6] = 32'b010000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [7] = 32'b010000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [8] = 32'b010000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [9] = 32'b010000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [10] = 32'b010000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [11] = 32'b010000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [12] = 32'b010000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [13] = 32'b010000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [14] = 32'b010000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [15] = 32'b010000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [16] = 32'b010000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [17] = 32'b010000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [18] = 32'b010000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [19] = 32'b010000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [20] = 32'b010000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [21] = 32'b010000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [22] = 32'b010000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [23] = 32'b010000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [24] = 32'b010000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [25] = 32'b010000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [26] = 32'b010000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [27] = 32'b010000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [28] = 32'b010000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [29] = 32'b010000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [30] = 32'b010000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r135 [31] = 32'b010000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [0] = 32'b010001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [1] = 32'b010001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [2] = 32'b010001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [3] = 32'b010001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [4] = 32'b010001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [5] = 32'b010001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [6] = 32'b010001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [7] = 32'b010001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [8] = 32'b010001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [9] = 32'b010001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [10] = 32'b010001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [11] = 32'b010001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [12] = 32'b010001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [13] = 32'b010001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [14] = 32'b010001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [15] = 32'b010001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [16] = 32'b010001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [17] = 32'b010001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [18] = 32'b010001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [19] = 32'b010001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [20] = 32'b010001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [21] = 32'b010001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [22] = 32'b010001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [23] = 32'b010001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [24] = 32'b010001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [25] = 32'b010001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [26] = 32'b010001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [27] = 32'b010001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [28] = 32'b010001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [29] = 32'b010001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [30] = 32'b010001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r134 [31] = 32'b010001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [0] = 32'b010001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [1] = 32'b010001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [2] = 32'b010001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [3] = 32'b010001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [4] = 32'b010001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [5] = 32'b010001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [6] = 32'b010001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [7] = 32'b010001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [8] = 32'b010001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [9] = 32'b010001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [10] = 32'b010001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [11] = 32'b010001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [12] = 32'b010001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [13] = 32'b010001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [14] = 32'b010001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [15] = 32'b010001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [16] = 32'b010001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [17] = 32'b010001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [18] = 32'b010001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [19] = 32'b010001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [20] = 32'b010001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [21] = 32'b010001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [22] = 32'b010001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [23] = 32'b010001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [24] = 32'b010001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [25] = 32'b010001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [26] = 32'b010001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [27] = 32'b010001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [28] = 32'b010001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [29] = 32'b010001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [30] = 32'b010001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r135 [31] = 32'b010001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [0] = 32'b010010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [1] = 32'b010010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [2] = 32'b010010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [3] = 32'b010010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [4] = 32'b010010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [5] = 32'b010010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [6] = 32'b010010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [7] = 32'b010010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [8] = 32'b010010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [9] = 32'b010010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [10] = 32'b010010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [11] = 32'b010010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [12] = 32'b010010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [13] = 32'b010010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [14] = 32'b010010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [15] = 32'b010010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [16] = 32'b010010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [17] = 32'b010010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [18] = 32'b010010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [19] = 32'b010010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [20] = 32'b010010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [21] = 32'b010010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [22] = 32'b010010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [23] = 32'b010010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [24] = 32'b010010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [25] = 32'b010010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [26] = 32'b010010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [27] = 32'b010010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [28] = 32'b010010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [29] = 32'b010010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [30] = 32'b010010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r134 [31] = 32'b010010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [0] = 32'b010010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [1] = 32'b010010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [2] = 32'b010010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [3] = 32'b010010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [4] = 32'b010010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [5] = 32'b010010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [6] = 32'b010010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [7] = 32'b010010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [8] = 32'b010010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [9] = 32'b010010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [10] = 32'b010010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [11] = 32'b010010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [12] = 32'b010010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [13] = 32'b010010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [14] = 32'b010010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [15] = 32'b010010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [16] = 32'b010010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [17] = 32'b010010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [18] = 32'b010010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [19] = 32'b010010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [20] = 32'b010010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [21] = 32'b010010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [22] = 32'b010010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [23] = 32'b010010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [24] = 32'b010010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [25] = 32'b010010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [26] = 32'b010010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [27] = 32'b010010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [28] = 32'b010010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [29] = 32'b010010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [30] = 32'b010010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r135 [31] = 32'b010010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [0] = 32'b010011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [1] = 32'b010011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [2] = 32'b010011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [3] = 32'b010011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [4] = 32'b010011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [5] = 32'b010011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [6] = 32'b010011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [7] = 32'b010011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [8] = 32'b010011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [9] = 32'b010011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [10] = 32'b010011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [11] = 32'b010011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [12] = 32'b010011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [13] = 32'b010011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [14] = 32'b010011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [15] = 32'b010011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [16] = 32'b010011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [17] = 32'b010011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [18] = 32'b010011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [19] = 32'b010011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [20] = 32'b010011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [21] = 32'b010011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [22] = 32'b010011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [23] = 32'b010011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [24] = 32'b010011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [25] = 32'b010011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [26] = 32'b010011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [27] = 32'b010011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [28] = 32'b010011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [29] = 32'b010011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [30] = 32'b010011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r134 [31] = 32'b010011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [0] = 32'b010011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [1] = 32'b010011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [2] = 32'b010011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [3] = 32'b010011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [4] = 32'b010011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [5] = 32'b010011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [6] = 32'b010011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [7] = 32'b010011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [8] = 32'b010011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [9] = 32'b010011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [10] = 32'b010011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [11] = 32'b010011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [12] = 32'b010011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [13] = 32'b010011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [14] = 32'b010011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [15] = 32'b010011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [16] = 32'b010011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [17] = 32'b010011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [18] = 32'b010011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [19] = 32'b010011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [20] = 32'b010011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [21] = 32'b010011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [22] = 32'b010011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [23] = 32'b010011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [24] = 32'b010011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [25] = 32'b010011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [26] = 32'b010011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [27] = 32'b010011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [28] = 32'b010011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [29] = 32'b010011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [30] = 32'b010011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r135 [31] = 32'b010011_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [0] = 32'b010100_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [1] = 32'b010100_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [2] = 32'b010100_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [3] = 32'b010100_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [4] = 32'b010100_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [5] = 32'b010100_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [6] = 32'b010100_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [7] = 32'b010100_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [8] = 32'b010100_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [9] = 32'b010100_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [10] = 32'b010100_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [11] = 32'b010100_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [12] = 32'b010100_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [13] = 32'b010100_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [14] = 32'b010100_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [15] = 32'b010100_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [16] = 32'b010100_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [17] = 32'b010100_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [18] = 32'b010100_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [19] = 32'b010100_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [20] = 32'b010100_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [21] = 32'b010100_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [22] = 32'b010100_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [23] = 32'b010100_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [24] = 32'b010100_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [25] = 32'b010100_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [26] = 32'b010100_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [27] = 32'b010100_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [28] = 32'b010100_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [29] = 32'b010100_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [30] = 32'b010100_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r134 [31] = 32'b010100_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [0] = 32'b010100_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [1] = 32'b010100_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [2] = 32'b010100_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [3] = 32'b010100_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [4] = 32'b010100_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [5] = 32'b010100_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [6] = 32'b010100_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [7] = 32'b010100_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [8] = 32'b010100_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [9] = 32'b010100_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [10] = 32'b010100_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [11] = 32'b010100_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [12] = 32'b010100_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [13] = 32'b010100_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [14] = 32'b010100_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [15] = 32'b010100_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [16] = 32'b010100_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [17] = 32'b010100_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [18] = 32'b010100_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [19] = 32'b010100_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [20] = 32'b010100_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [21] = 32'b010100_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [22] = 32'b010100_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [23] = 32'b010100_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [24] = 32'b010100_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [25] = 32'b010100_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [26] = 32'b010100_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [27] = 32'b010100_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [28] = 32'b010100_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [29] = 32'b010100_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [30] = 32'b010100_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r135 [31] = 32'b010100_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [0] = 32'b010101_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [1] = 32'b010101_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [2] = 32'b010101_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [3] = 32'b010101_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [4] = 32'b010101_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [5] = 32'b010101_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [6] = 32'b010101_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [7] = 32'b010101_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [8] = 32'b010101_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [9] = 32'b010101_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [10] = 32'b010101_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [11] = 32'b010101_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [12] = 32'b010101_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [13] = 32'b010101_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [14] = 32'b010101_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [15] = 32'b010101_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [16] = 32'b010101_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [17] = 32'b010101_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [18] = 32'b010101_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [19] = 32'b010101_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [20] = 32'b010101_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [21] = 32'b010101_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [22] = 32'b010101_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [23] = 32'b010101_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [24] = 32'b010101_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [25] = 32'b010101_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [26] = 32'b010101_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [27] = 32'b010101_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [28] = 32'b010101_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [29] = 32'b010101_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [30] = 32'b010101_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r134 [31] = 32'b010101_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [0] = 32'b010101_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [1] = 32'b010101_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [2] = 32'b010101_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [3] = 32'b010101_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [4] = 32'b010101_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [5] = 32'b010101_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [6] = 32'b010101_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [7] = 32'b010101_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [8] = 32'b010101_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [9] = 32'b010101_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [10] = 32'b010101_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [11] = 32'b010101_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [12] = 32'b010101_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [13] = 32'b010101_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [14] = 32'b010101_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [15] = 32'b010101_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [16] = 32'b010101_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [17] = 32'b010101_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [18] = 32'b010101_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [19] = 32'b010101_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [20] = 32'b010101_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [21] = 32'b010101_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [22] = 32'b010101_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [23] = 32'b010101_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [24] = 32'b010101_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [25] = 32'b010101_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [26] = 32'b010101_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [27] = 32'b010101_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [28] = 32'b010101_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [29] = 32'b010101_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [30] = 32'b010101_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r135 [31] = 32'b010101_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [0] = 32'b010110_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [1] = 32'b010110_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [2] = 32'b010110_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [3] = 32'b010110_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [4] = 32'b010110_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [5] = 32'b010110_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [6] = 32'b010110_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [7] = 32'b010110_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [8] = 32'b010110_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [9] = 32'b010110_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [10] = 32'b010110_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [11] = 32'b010110_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [12] = 32'b010110_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [13] = 32'b010110_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [14] = 32'b010110_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [15] = 32'b010110_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [16] = 32'b010110_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [17] = 32'b010110_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [18] = 32'b010110_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [19] = 32'b010110_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [20] = 32'b010110_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [21] = 32'b010110_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [22] = 32'b010110_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [23] = 32'b010110_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [24] = 32'b010110_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [25] = 32'b010110_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [26] = 32'b010110_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [27] = 32'b010110_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [28] = 32'b010110_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [29] = 32'b010110_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [30] = 32'b010110_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r134 [31] = 32'b010110_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [0] = 32'b010110_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [1] = 32'b010110_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [2] = 32'b010110_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [3] = 32'b010110_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [4] = 32'b010110_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [5] = 32'b010110_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [6] = 32'b010110_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [7] = 32'b010110_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [8] = 32'b010110_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [9] = 32'b010110_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [10] = 32'b010110_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [11] = 32'b010110_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [12] = 32'b010110_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [13] = 32'b010110_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [14] = 32'b010110_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [15] = 32'b010110_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [16] = 32'b010110_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [17] = 32'b010110_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [18] = 32'b010110_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [19] = 32'b010110_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [20] = 32'b010110_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [21] = 32'b010110_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [22] = 32'b010110_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [23] = 32'b010110_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [24] = 32'b010110_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [25] = 32'b010110_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [26] = 32'b010110_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [27] = 32'b010110_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [28] = 32'b010110_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [29] = 32'b010110_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [30] = 32'b010110_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r135 [31] = 32'b010110_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [0] = 32'b010111_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [1] = 32'b010111_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [2] = 32'b010111_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [3] = 32'b010111_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [4] = 32'b010111_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [5] = 32'b010111_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [6] = 32'b010111_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [7] = 32'b010111_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [8] = 32'b010111_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [9] = 32'b010111_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [10] = 32'b010111_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [11] = 32'b010111_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [12] = 32'b010111_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [13] = 32'b010111_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [14] = 32'b010111_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [15] = 32'b010111_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [16] = 32'b010111_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [17] = 32'b010111_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [18] = 32'b010111_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [19] = 32'b010111_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [20] = 32'b010111_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [21] = 32'b010111_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [22] = 32'b010111_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [23] = 32'b010111_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [24] = 32'b010111_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [25] = 32'b010111_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [26] = 32'b010111_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [27] = 32'b010111_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [28] = 32'b010111_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [29] = 32'b010111_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [30] = 32'b010111_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r134 [31] = 32'b010111_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [0] = 32'b010111_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [1] = 32'b010111_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [2] = 32'b010111_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [3] = 32'b010111_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [4] = 32'b010111_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [5] = 32'b010111_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [6] = 32'b010111_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [7] = 32'b010111_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [8] = 32'b010111_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [9] = 32'b010111_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [10] = 32'b010111_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [11] = 32'b010111_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [12] = 32'b010111_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [13] = 32'b010111_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [14] = 32'b010111_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [15] = 32'b010111_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [16] = 32'b010111_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [17] = 32'b010111_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [18] = 32'b010111_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [19] = 32'b010111_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [20] = 32'b010111_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [21] = 32'b010111_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [22] = 32'b010111_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [23] = 32'b010111_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [24] = 32'b010111_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [25] = 32'b010111_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [26] = 32'b010111_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [27] = 32'b010111_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [28] = 32'b010111_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [29] = 32'b010111_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [30] = 32'b010111_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r135 [31] = 32'b010111_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [0] = 32'b011000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [1] = 32'b011000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [2] = 32'b011000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [3] = 32'b011000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [4] = 32'b011000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [5] = 32'b011000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [6] = 32'b011000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [7] = 32'b011000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [8] = 32'b011000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [9] = 32'b011000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [10] = 32'b011000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [11] = 32'b011000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [12] = 32'b011000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [13] = 32'b011000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [14] = 32'b011000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [15] = 32'b011000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [16] = 32'b011000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [17] = 32'b011000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [18] = 32'b011000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [19] = 32'b011000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [20] = 32'b011000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [21] = 32'b011000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [22] = 32'b011000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [23] = 32'b011000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [24] = 32'b011000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [25] = 32'b011000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [26] = 32'b011000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [27] = 32'b011000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [28] = 32'b011000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [29] = 32'b011000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [30] = 32'b011000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r134 [31] = 32'b011000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [0] = 32'b011000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [1] = 32'b011000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [2] = 32'b011000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [3] = 32'b011000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [4] = 32'b011000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [5] = 32'b011000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [6] = 32'b011000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [7] = 32'b011000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [8] = 32'b011000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [9] = 32'b011000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [10] = 32'b011000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [11] = 32'b011000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [12] = 32'b011000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [13] = 32'b011000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [14] = 32'b011000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [15] = 32'b011000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [16] = 32'b011000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [17] = 32'b011000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [18] = 32'b011000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [19] = 32'b011000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [20] = 32'b011000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [21] = 32'b011000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [22] = 32'b011000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [23] = 32'b011000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [24] = 32'b011000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [25] = 32'b011000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [26] = 32'b011000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [27] = 32'b011000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [28] = 32'b011000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [29] = 32'b011000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [30] = 32'b011000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r135 [31] = 32'b011000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [0] = 32'b011001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [1] = 32'b011001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [2] = 32'b011001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [3] = 32'b011001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [4] = 32'b011001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [5] = 32'b011001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [6] = 32'b011001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [7] = 32'b011001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [8] = 32'b011001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [9] = 32'b011001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [10] = 32'b011001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [11] = 32'b011001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [12] = 32'b011001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [13] = 32'b011001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [14] = 32'b011001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [15] = 32'b011001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [16] = 32'b011001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [17] = 32'b011001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [18] = 32'b011001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [19] = 32'b011001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [20] = 32'b011001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [21] = 32'b011001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [22] = 32'b011001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [23] = 32'b011001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [24] = 32'b011001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [25] = 32'b011001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [26] = 32'b011001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [27] = 32'b011001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [28] = 32'b011001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [29] = 32'b011001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [30] = 32'b011001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r134 [31] = 32'b011001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [0] = 32'b011001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [1] = 32'b011001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [2] = 32'b011001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [3] = 32'b011001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [4] = 32'b011001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [5] = 32'b011001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [6] = 32'b011001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [7] = 32'b011001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [8] = 32'b011001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [9] = 32'b011001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [10] = 32'b011001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [11] = 32'b011001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [12] = 32'b011001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [13] = 32'b011001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [14] = 32'b011001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [15] = 32'b011001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [16] = 32'b011001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [17] = 32'b011001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [18] = 32'b011001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [19] = 32'b011001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [20] = 32'b011001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [21] = 32'b011001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [22] = 32'b011001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [23] = 32'b011001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [24] = 32'b011001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [25] = 32'b011001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [26] = 32'b011001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [27] = 32'b011001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [28] = 32'b011001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [29] = 32'b011001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [30] = 32'b011001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r135 [31] = 32'b011001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [0] = 32'b011010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [1] = 32'b011010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [2] = 32'b011010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [3] = 32'b011010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [4] = 32'b011010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [5] = 32'b011010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [6] = 32'b011010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [7] = 32'b011010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [8] = 32'b011010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [9] = 32'b011010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [10] = 32'b011010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [11] = 32'b011010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [12] = 32'b011010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [13] = 32'b011010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [14] = 32'b011010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [15] = 32'b011010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [16] = 32'b011010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [17] = 32'b011010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [18] = 32'b011010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [19] = 32'b011010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [20] = 32'b011010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [21] = 32'b011010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [22] = 32'b011010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [23] = 32'b011010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [24] = 32'b011010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [25] = 32'b011010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [26] = 32'b011010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [27] = 32'b011010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [28] = 32'b011010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [29] = 32'b011010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [30] = 32'b011010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r134 [31] = 32'b011010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [0] = 32'b011010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [1] = 32'b011010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [2] = 32'b011010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [3] = 32'b011010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [4] = 32'b011010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [5] = 32'b011010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [6] = 32'b011010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [7] = 32'b011010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [8] = 32'b011010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [9] = 32'b011010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [10] = 32'b011010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [11] = 32'b011010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [12] = 32'b011010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [13] = 32'b011010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [14] = 32'b011010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [15] = 32'b011010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [16] = 32'b011010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [17] = 32'b011010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [18] = 32'b011010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [19] = 32'b011010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [20] = 32'b011010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [21] = 32'b011010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [22] = 32'b011010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [23] = 32'b011010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [24] = 32'b011010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [25] = 32'b011010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [26] = 32'b011010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [27] = 32'b011010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [28] = 32'b011010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [29] = 32'b011010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [30] = 32'b011010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r135 [31] = 32'b011010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [0] = 32'b011011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [1] = 32'b011011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [2] = 32'b011011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [3] = 32'b011011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [4] = 32'b011011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [5] = 32'b011011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [6] = 32'b011011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [7] = 32'b011011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [8] = 32'b011011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [9] = 32'b011011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [10] = 32'b011011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [11] = 32'b011011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [12] = 32'b011011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [13] = 32'b011011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [14] = 32'b011011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [15] = 32'b011011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [16] = 32'b011011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [17] = 32'b011011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [18] = 32'b011011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [19] = 32'b011011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [20] = 32'b011011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [21] = 32'b011011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [22] = 32'b011011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [23] = 32'b011011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [24] = 32'b011011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [25] = 32'b011011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [26] = 32'b011011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [27] = 32'b011011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [28] = 32'b011011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [29] = 32'b011011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [30] = 32'b011011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r134 [31] = 32'b011011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [0] = 32'b011011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [1] = 32'b011011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [2] = 32'b011011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [3] = 32'b011011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [4] = 32'b011011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [5] = 32'b011011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [6] = 32'b011011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [7] = 32'b011011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [8] = 32'b011011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [9] = 32'b011011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [10] = 32'b011011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [11] = 32'b011011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [12] = 32'b011011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [13] = 32'b011011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [14] = 32'b011011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [15] = 32'b011011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [16] = 32'b011011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [17] = 32'b011011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [18] = 32'b011011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [19] = 32'b011011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [20] = 32'b011011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [21] = 32'b011011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [22] = 32'b011011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [23] = 32'b011011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [24] = 32'b011011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [25] = 32'b011011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [26] = 32'b011011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [27] = 32'b011011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [28] = 32'b011011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [29] = 32'b011011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [30] = 32'b011011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r135 [31] = 32'b011011_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [0] = 32'b011100_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [1] = 32'b011100_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [2] = 32'b011100_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [3] = 32'b011100_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [4] = 32'b011100_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [5] = 32'b011100_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [6] = 32'b011100_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [7] = 32'b011100_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [8] = 32'b011100_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [9] = 32'b011100_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [10] = 32'b011100_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [11] = 32'b011100_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [12] = 32'b011100_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [13] = 32'b011100_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [14] = 32'b011100_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [15] = 32'b011100_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [16] = 32'b011100_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [17] = 32'b011100_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [18] = 32'b011100_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [19] = 32'b011100_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [20] = 32'b011100_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [21] = 32'b011100_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [22] = 32'b011100_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [23] = 32'b011100_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [24] = 32'b011100_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [25] = 32'b011100_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [26] = 32'b011100_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [27] = 32'b011100_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [28] = 32'b011100_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [29] = 32'b011100_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [30] = 32'b011100_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r134 [31] = 32'b011100_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [0] = 32'b011100_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [1] = 32'b011100_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [2] = 32'b011100_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [3] = 32'b011100_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [4] = 32'b011100_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [5] = 32'b011100_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [6] = 32'b011100_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [7] = 32'b011100_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [8] = 32'b011100_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [9] = 32'b011100_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [10] = 32'b011100_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [11] = 32'b011100_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [12] = 32'b011100_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [13] = 32'b011100_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [14] = 32'b011100_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [15] = 32'b011100_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [16] = 32'b011100_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [17] = 32'b011100_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [18] = 32'b011100_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [19] = 32'b011100_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [20] = 32'b011100_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [21] = 32'b011100_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [22] = 32'b011100_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [23] = 32'b011100_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [24] = 32'b011100_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [25] = 32'b011100_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [26] = 32'b011100_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [27] = 32'b011100_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [28] = 32'b011100_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [29] = 32'b011100_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [30] = 32'b011100_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r135 [31] = 32'b011100_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [0] = 32'b011101_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [1] = 32'b011101_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [2] = 32'b011101_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [3] = 32'b011101_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [4] = 32'b011101_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [5] = 32'b011101_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [6] = 32'b011101_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [7] = 32'b011101_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [8] = 32'b011101_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [9] = 32'b011101_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [10] = 32'b011101_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [11] = 32'b011101_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [12] = 32'b011101_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [13] = 32'b011101_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [14] = 32'b011101_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [15] = 32'b011101_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [16] = 32'b011101_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [17] = 32'b011101_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [18] = 32'b011101_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [19] = 32'b011101_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [20] = 32'b011101_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [21] = 32'b011101_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [22] = 32'b011101_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [23] = 32'b011101_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [24] = 32'b011101_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [25] = 32'b011101_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [26] = 32'b011101_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [27] = 32'b011101_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [28] = 32'b011101_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [29] = 32'b011101_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [30] = 32'b011101_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r134 [31] = 32'b011101_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [0] = 32'b011101_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [1] = 32'b011101_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [2] = 32'b011101_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [3] = 32'b011101_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [4] = 32'b011101_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [5] = 32'b011101_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [6] = 32'b011101_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [7] = 32'b011101_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [8] = 32'b011101_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [9] = 32'b011101_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [10] = 32'b011101_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [11] = 32'b011101_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [12] = 32'b011101_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [13] = 32'b011101_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [14] = 32'b011101_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [15] = 32'b011101_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [16] = 32'b011101_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [17] = 32'b011101_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [18] = 32'b011101_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [19] = 32'b011101_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [20] = 32'b011101_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [21] = 32'b011101_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [22] = 32'b011101_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [23] = 32'b011101_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [24] = 32'b011101_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [25] = 32'b011101_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [26] = 32'b011101_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [27] = 32'b011101_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [28] = 32'b011101_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [29] = 32'b011101_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [30] = 32'b011101_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r135 [31] = 32'b011101_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [0] = 32'b011110_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [1] = 32'b011110_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [2] = 32'b011110_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [3] = 32'b011110_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [4] = 32'b011110_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [5] = 32'b011110_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [6] = 32'b011110_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [7] = 32'b011110_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [8] = 32'b011110_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [9] = 32'b011110_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [10] = 32'b011110_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [11] = 32'b011110_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [12] = 32'b011110_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [13] = 32'b011110_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [14] = 32'b011110_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [15] = 32'b011110_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [16] = 32'b011110_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [17] = 32'b011110_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [18] = 32'b011110_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [19] = 32'b011110_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [20] = 32'b011110_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [21] = 32'b011110_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [22] = 32'b011110_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [23] = 32'b011110_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [24] = 32'b011110_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [25] = 32'b011110_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [26] = 32'b011110_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [27] = 32'b011110_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [28] = 32'b011110_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [29] = 32'b011110_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [30] = 32'b011110_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r134 [31] = 32'b011110_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [0] = 32'b011110_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [1] = 32'b011110_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [2] = 32'b011110_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [3] = 32'b011110_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [4] = 32'b011110_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [5] = 32'b011110_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [6] = 32'b011110_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [7] = 32'b011110_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [8] = 32'b011110_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [9] = 32'b011110_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [10] = 32'b011110_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [11] = 32'b011110_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [12] = 32'b011110_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [13] = 32'b011110_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [14] = 32'b011110_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [15] = 32'b011110_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [16] = 32'b011110_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [17] = 32'b011110_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [18] = 32'b011110_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [19] = 32'b011110_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [20] = 32'b011110_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [21] = 32'b011110_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [22] = 32'b011110_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [23] = 32'b011110_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [24] = 32'b011110_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [25] = 32'b011110_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [26] = 32'b011110_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [27] = 32'b011110_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [28] = 32'b011110_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [29] = 32'b011110_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [30] = 32'b011110_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r135 [31] = 32'b011110_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [0] = 32'b011111_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [1] = 32'b011111_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [2] = 32'b011111_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [3] = 32'b011111_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [4] = 32'b011111_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [5] = 32'b011111_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [6] = 32'b011111_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [7] = 32'b011111_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [8] = 32'b011111_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [9] = 32'b011111_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [10] = 32'b011111_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [11] = 32'b011111_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [12] = 32'b011111_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [13] = 32'b011111_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [14] = 32'b011111_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [15] = 32'b011111_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [16] = 32'b011111_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [17] = 32'b011111_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [18] = 32'b011111_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [19] = 32'b011111_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [20] = 32'b011111_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [21] = 32'b011111_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [22] = 32'b011111_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [23] = 32'b011111_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [24] = 32'b011111_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [25] = 32'b011111_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [26] = 32'b011111_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [27] = 32'b011111_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [28] = 32'b011111_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [29] = 32'b011111_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [30] = 32'b011111_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r134 [31] = 32'b011111_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [0] = 32'b011111_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [1] = 32'b011111_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [2] = 32'b011111_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [3] = 32'b011111_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [4] = 32'b011111_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [5] = 32'b011111_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [6] = 32'b011111_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [7] = 32'b011111_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [8] = 32'b011111_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [9] = 32'b011111_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [10] = 32'b011111_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [11] = 32'b011111_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [12] = 32'b011111_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [13] = 32'b011111_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [14] = 32'b011111_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [15] = 32'b011111_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [16] = 32'b011111_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [17] = 32'b011111_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [18] = 32'b011111_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [19] = 32'b011111_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [20] = 32'b011111_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [21] = 32'b011111_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [22] = 32'b011111_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [23] = 32'b011111_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [24] = 32'b011111_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [25] = 32'b011111_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [26] = 32'b011111_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [27] = 32'b011111_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [28] = 32'b011111_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [29] = 32'b011111_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [30] = 32'b011111_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r135 [31] = 32'b011111_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [0] = 32'b100000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [1] = 32'b100000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [2] = 32'b100000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [3] = 32'b100000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [4] = 32'b100000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [5] = 32'b100000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [6] = 32'b100000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [7] = 32'b100000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [8] = 32'b100000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [9] = 32'b100000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [10] = 32'b100000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [11] = 32'b100000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [12] = 32'b100000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [13] = 32'b100000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [14] = 32'b100000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [15] = 32'b100000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [16] = 32'b100000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [17] = 32'b100000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [18] = 32'b100000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [19] = 32'b100000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [20] = 32'b100000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [21] = 32'b100000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [22] = 32'b100000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [23] = 32'b100000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [24] = 32'b100000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [25] = 32'b100000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [26] = 32'b100000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [27] = 32'b100000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [28] = 32'b100000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [29] = 32'b100000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [30] = 32'b100000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r134 [31] = 32'b100000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [0] = 32'b100000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [1] = 32'b100000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [2] = 32'b100000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [3] = 32'b100000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [4] = 32'b100000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [5] = 32'b100000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [6] = 32'b100000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [7] = 32'b100000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [8] = 32'b100000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [9] = 32'b100000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [10] = 32'b100000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [11] = 32'b100000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [12] = 32'b100000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [13] = 32'b100000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [14] = 32'b100000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [15] = 32'b100000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [16] = 32'b100000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [17] = 32'b100000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [18] = 32'b100000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [19] = 32'b100000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [20] = 32'b100000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [21] = 32'b100000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [22] = 32'b100000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [23] = 32'b100000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [24] = 32'b100000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [25] = 32'b100000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [26] = 32'b100000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [27] = 32'b100000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [28] = 32'b100000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [29] = 32'b100000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [30] = 32'b100000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r135 [31] = 32'b100000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [0] = 32'b100001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [1] = 32'b100001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [2] = 32'b100001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [3] = 32'b100001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [4] = 32'b100001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [5] = 32'b100001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [6] = 32'b100001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [7] = 32'b100001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [8] = 32'b100001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [9] = 32'b100001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [10] = 32'b100001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [11] = 32'b100001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [12] = 32'b100001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [13] = 32'b100001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [14] = 32'b100001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [15] = 32'b100001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [16] = 32'b100001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [17] = 32'b100001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [18] = 32'b100001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [19] = 32'b100001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [20] = 32'b100001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [21] = 32'b100001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [22] = 32'b100001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [23] = 32'b100001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [24] = 32'b100001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [25] = 32'b100001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [26] = 32'b100001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [27] = 32'b100001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [28] = 32'b100001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [29] = 32'b100001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [30] = 32'b100001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r134 [31] = 32'b100001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [0] = 32'b100001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [1] = 32'b100001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [2] = 32'b100001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [3] = 32'b100001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [4] = 32'b100001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [5] = 32'b100001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [6] = 32'b100001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [7] = 32'b100001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [8] = 32'b100001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [9] = 32'b100001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [10] = 32'b100001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [11] = 32'b100001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [12] = 32'b100001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [13] = 32'b100001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [14] = 32'b100001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [15] = 32'b100001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [16] = 32'b100001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [17] = 32'b100001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [18] = 32'b100001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [19] = 32'b100001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [20] = 32'b100001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [21] = 32'b100001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [22] = 32'b100001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [23] = 32'b100001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [24] = 32'b100001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [25] = 32'b100001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [26] = 32'b100001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [27] = 32'b100001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [28] = 32'b100001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [29] = 32'b100001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [30] = 32'b100001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r135 [31] = 32'b100001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [0] = 32'b100010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [1] = 32'b100010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [2] = 32'b100010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [3] = 32'b100010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [4] = 32'b100010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [5] = 32'b100010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [6] = 32'b100010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [7] = 32'b100010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [8] = 32'b100010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [9] = 32'b100010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [10] = 32'b100010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [11] = 32'b100010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [12] = 32'b100010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [13] = 32'b100010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [14] = 32'b100010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [15] = 32'b100010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [16] = 32'b100010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [17] = 32'b100010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [18] = 32'b100010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [19] = 32'b100010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [20] = 32'b100010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [21] = 32'b100010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [22] = 32'b100010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [23] = 32'b100010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [24] = 32'b100010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [25] = 32'b100010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [26] = 32'b100010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [27] = 32'b100010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [28] = 32'b100010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [29] = 32'b100010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [30] = 32'b100010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r134 [31] = 32'b100010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [0] = 32'b100010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [1] = 32'b100010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [2] = 32'b100010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [3] = 32'b100010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [4] = 32'b100010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [5] = 32'b100010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [6] = 32'b100010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [7] = 32'b100010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [8] = 32'b100010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [9] = 32'b100010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [10] = 32'b100010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [11] = 32'b100010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [12] = 32'b100010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [13] = 32'b100010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [14] = 32'b100010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [15] = 32'b100010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [16] = 32'b100010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [17] = 32'b100010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [18] = 32'b100010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [19] = 32'b100010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [20] = 32'b100010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [21] = 32'b100010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [22] = 32'b100010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [23] = 32'b100010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [24] = 32'b100010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [25] = 32'b100010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [26] = 32'b100010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [27] = 32'b100010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [28] = 32'b100010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [29] = 32'b100010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [30] = 32'b100010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r135 [31] = 32'b100010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [0] = 32'b100011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [1] = 32'b100011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [2] = 32'b100011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [3] = 32'b100011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [4] = 32'b100011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [5] = 32'b100011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [6] = 32'b100011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [7] = 32'b100011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [8] = 32'b100011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [9] = 32'b100011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [10] = 32'b100011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [11] = 32'b100011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [12] = 32'b100011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [13] = 32'b100011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [14] = 32'b100011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [15] = 32'b100011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [16] = 32'b100011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [17] = 32'b100011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [18] = 32'b100011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [19] = 32'b100011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [20] = 32'b100011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [21] = 32'b100011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [22] = 32'b100011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [23] = 32'b100011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [24] = 32'b100011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [25] = 32'b100011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [26] = 32'b100011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [27] = 32'b100011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [28] = 32'b100011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [29] = 32'b100011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [30] = 32'b100011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r134 [31] = 32'b100011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [0] = 32'b100011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [1] = 32'b100011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [2] = 32'b100011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [3] = 32'b100011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [4] = 32'b100011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [5] = 32'b100011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [6] = 32'b100011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [7] = 32'b100011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [8] = 32'b100011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [9] = 32'b100011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [10] = 32'b100011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [11] = 32'b100011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [12] = 32'b100011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [13] = 32'b100011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [14] = 32'b100011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [15] = 32'b100011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [16] = 32'b100011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [17] = 32'b100011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [18] = 32'b100011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [19] = 32'b100011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [20] = 32'b100011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [21] = 32'b100011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [22] = 32'b100011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [23] = 32'b100011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [24] = 32'b100011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [25] = 32'b100011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [26] = 32'b100011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [27] = 32'b100011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [28] = 32'b100011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [29] = 32'b100011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [30] = 32'b100011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r135 [31] = 32'b100011_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [0] = 32'b100100_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [1] = 32'b100100_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [2] = 32'b100100_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [3] = 32'b100100_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [4] = 32'b100100_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [5] = 32'b100100_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [6] = 32'b100100_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [7] = 32'b100100_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [8] = 32'b100100_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [9] = 32'b100100_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [10] = 32'b100100_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [11] = 32'b100100_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [12] = 32'b100100_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [13] = 32'b100100_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [14] = 32'b100100_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [15] = 32'b100100_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [16] = 32'b100100_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [17] = 32'b100100_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [18] = 32'b100100_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [19] = 32'b100100_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [20] = 32'b100100_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [21] = 32'b100100_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [22] = 32'b100100_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [23] = 32'b100100_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [24] = 32'b100100_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [25] = 32'b100100_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [26] = 32'b100100_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [27] = 32'b100100_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [28] = 32'b100100_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [29] = 32'b100100_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [30] = 32'b100100_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r134 [31] = 32'b100100_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [0] = 32'b100100_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [1] = 32'b100100_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [2] = 32'b100100_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [3] = 32'b100100_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [4] = 32'b100100_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [5] = 32'b100100_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [6] = 32'b100100_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [7] = 32'b100100_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [8] = 32'b100100_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [9] = 32'b100100_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [10] = 32'b100100_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [11] = 32'b100100_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [12] = 32'b100100_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [13] = 32'b100100_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [14] = 32'b100100_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [15] = 32'b100100_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [16] = 32'b100100_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [17] = 32'b100100_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [18] = 32'b100100_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [19] = 32'b100100_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [20] = 32'b100100_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [21] = 32'b100100_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [22] = 32'b100100_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [23] = 32'b100100_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [24] = 32'b100100_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [25] = 32'b100100_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [26] = 32'b100100_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [27] = 32'b100100_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [28] = 32'b100100_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [29] = 32'b100100_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [30] = 32'b100100_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r135 [31] = 32'b100100_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [0] = 32'b100101_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [1] = 32'b100101_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [2] = 32'b100101_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [3] = 32'b100101_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [4] = 32'b100101_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [5] = 32'b100101_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [6] = 32'b100101_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [7] = 32'b100101_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [8] = 32'b100101_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [9] = 32'b100101_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [10] = 32'b100101_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [11] = 32'b100101_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [12] = 32'b100101_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [13] = 32'b100101_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [14] = 32'b100101_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [15] = 32'b100101_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [16] = 32'b100101_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [17] = 32'b100101_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [18] = 32'b100101_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [19] = 32'b100101_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [20] = 32'b100101_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [21] = 32'b100101_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [22] = 32'b100101_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [23] = 32'b100101_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [24] = 32'b100101_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [25] = 32'b100101_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [26] = 32'b100101_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [27] = 32'b100101_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [28] = 32'b100101_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [29] = 32'b100101_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [30] = 32'b100101_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r134 [31] = 32'b100101_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [0] = 32'b100101_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [1] = 32'b100101_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [2] = 32'b100101_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [3] = 32'b100101_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [4] = 32'b100101_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [5] = 32'b100101_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [6] = 32'b100101_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [7] = 32'b100101_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [8] = 32'b100101_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [9] = 32'b100101_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [10] = 32'b100101_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [11] = 32'b100101_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [12] = 32'b100101_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [13] = 32'b100101_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [14] = 32'b100101_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [15] = 32'b100101_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [16] = 32'b100101_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [17] = 32'b100101_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [18] = 32'b100101_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [19] = 32'b100101_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [20] = 32'b100101_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [21] = 32'b100101_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [22] = 32'b100101_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [23] = 32'b100101_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [24] = 32'b100101_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [25] = 32'b100101_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [26] = 32'b100101_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [27] = 32'b100101_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [28] = 32'b100101_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [29] = 32'b100101_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [30] = 32'b100101_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r135 [31] = 32'b100101_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [0] = 32'b100110_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [1] = 32'b100110_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [2] = 32'b100110_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [3] = 32'b100110_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [4] = 32'b100110_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [5] = 32'b100110_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [6] = 32'b100110_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [7] = 32'b100110_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [8] = 32'b100110_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [9] = 32'b100110_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [10] = 32'b100110_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [11] = 32'b100110_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [12] = 32'b100110_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [13] = 32'b100110_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [14] = 32'b100110_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [15] = 32'b100110_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [16] = 32'b100110_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [17] = 32'b100110_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [18] = 32'b100110_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [19] = 32'b100110_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [20] = 32'b100110_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [21] = 32'b100110_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [22] = 32'b100110_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [23] = 32'b100110_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [24] = 32'b100110_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [25] = 32'b100110_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [26] = 32'b100110_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [27] = 32'b100110_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [28] = 32'b100110_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [29] = 32'b100110_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [30] = 32'b100110_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r134 [31] = 32'b100110_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [0] = 32'b100110_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [1] = 32'b100110_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [2] = 32'b100110_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [3] = 32'b100110_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [4] = 32'b100110_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [5] = 32'b100110_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [6] = 32'b100110_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [7] = 32'b100110_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [8] = 32'b100110_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [9] = 32'b100110_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [10] = 32'b100110_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [11] = 32'b100110_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [12] = 32'b100110_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [13] = 32'b100110_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [14] = 32'b100110_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [15] = 32'b100110_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [16] = 32'b100110_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [17] = 32'b100110_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [18] = 32'b100110_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [19] = 32'b100110_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [20] = 32'b100110_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [21] = 32'b100110_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [22] = 32'b100110_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [23] = 32'b100110_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [24] = 32'b100110_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [25] = 32'b100110_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [26] = 32'b100110_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [27] = 32'b100110_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [28] = 32'b100110_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [29] = 32'b100110_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [30] = 32'b100110_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r135 [31] = 32'b100110_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [0] = 32'b100111_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [1] = 32'b100111_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [2] = 32'b100111_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [3] = 32'b100111_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [4] = 32'b100111_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [5] = 32'b100111_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [6] = 32'b100111_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [7] = 32'b100111_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [8] = 32'b100111_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [9] = 32'b100111_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [10] = 32'b100111_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [11] = 32'b100111_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [12] = 32'b100111_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [13] = 32'b100111_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [14] = 32'b100111_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [15] = 32'b100111_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [16] = 32'b100111_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [17] = 32'b100111_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [18] = 32'b100111_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [19] = 32'b100111_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [20] = 32'b100111_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [21] = 32'b100111_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [22] = 32'b100111_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [23] = 32'b100111_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [24] = 32'b100111_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [25] = 32'b100111_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [26] = 32'b100111_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [27] = 32'b100111_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [28] = 32'b100111_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [29] = 32'b100111_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [30] = 32'b100111_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r134 [31] = 32'b100111_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [0] = 32'b100111_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [1] = 32'b100111_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [2] = 32'b100111_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [3] = 32'b100111_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [4] = 32'b100111_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [5] = 32'b100111_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [6] = 32'b100111_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [7] = 32'b100111_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [8] = 32'b100111_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [9] = 32'b100111_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [10] = 32'b100111_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [11] = 32'b100111_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [12] = 32'b100111_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [13] = 32'b100111_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [14] = 32'b100111_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [15] = 32'b100111_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [16] = 32'b100111_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [17] = 32'b100111_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [18] = 32'b100111_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [19] = 32'b100111_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [20] = 32'b100111_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [21] = 32'b100111_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [22] = 32'b100111_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [23] = 32'b100111_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [24] = 32'b100111_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [25] = 32'b100111_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [26] = 32'b100111_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [27] = 32'b100111_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [28] = 32'b100111_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [29] = 32'b100111_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [30] = 32'b100111_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r135 [31] = 32'b100111_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [0] = 32'b101000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [1] = 32'b101000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [2] = 32'b101000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [3] = 32'b101000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [4] = 32'b101000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [5] = 32'b101000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [6] = 32'b101000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [7] = 32'b101000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [8] = 32'b101000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [9] = 32'b101000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [10] = 32'b101000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [11] = 32'b101000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [12] = 32'b101000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [13] = 32'b101000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [14] = 32'b101000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [15] = 32'b101000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [16] = 32'b101000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [17] = 32'b101000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [18] = 32'b101000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [19] = 32'b101000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [20] = 32'b101000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [21] = 32'b101000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [22] = 32'b101000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [23] = 32'b101000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [24] = 32'b101000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [25] = 32'b101000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [26] = 32'b101000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [27] = 32'b101000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [28] = 32'b101000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [29] = 32'b101000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [30] = 32'b101000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r134 [31] = 32'b101000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [0] = 32'b101000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [1] = 32'b101000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [2] = 32'b101000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [3] = 32'b101000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [4] = 32'b101000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [5] = 32'b101000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [6] = 32'b101000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [7] = 32'b101000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [8] = 32'b101000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [9] = 32'b101000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [10] = 32'b101000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [11] = 32'b101000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [12] = 32'b101000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [13] = 32'b101000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [14] = 32'b101000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [15] = 32'b101000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [16] = 32'b101000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [17] = 32'b101000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [18] = 32'b101000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [19] = 32'b101000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [20] = 32'b101000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [21] = 32'b101000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [22] = 32'b101000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [23] = 32'b101000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [24] = 32'b101000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [25] = 32'b101000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [26] = 32'b101000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [27] = 32'b101000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [28] = 32'b101000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [29] = 32'b101000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [30] = 32'b101000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r135 [31] = 32'b101000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [0] = 32'b101001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [1] = 32'b101001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [2] = 32'b101001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [3] = 32'b101001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [4] = 32'b101001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [5] = 32'b101001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [6] = 32'b101001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [7] = 32'b101001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [8] = 32'b101001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [9] = 32'b101001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [10] = 32'b101001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [11] = 32'b101001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [12] = 32'b101001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [13] = 32'b101001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [14] = 32'b101001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [15] = 32'b101001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [16] = 32'b101001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [17] = 32'b101001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [18] = 32'b101001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [19] = 32'b101001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [20] = 32'b101001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [21] = 32'b101001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [22] = 32'b101001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [23] = 32'b101001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [24] = 32'b101001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [25] = 32'b101001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [26] = 32'b101001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [27] = 32'b101001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [28] = 32'b101001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [29] = 32'b101001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [30] = 32'b101001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r134 [31] = 32'b101001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [0] = 32'b101001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [1] = 32'b101001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [2] = 32'b101001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [3] = 32'b101001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [4] = 32'b101001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [5] = 32'b101001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [6] = 32'b101001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [7] = 32'b101001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [8] = 32'b101001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [9] = 32'b101001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [10] = 32'b101001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [11] = 32'b101001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [12] = 32'b101001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [13] = 32'b101001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [14] = 32'b101001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [15] = 32'b101001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [16] = 32'b101001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [17] = 32'b101001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [18] = 32'b101001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [19] = 32'b101001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [20] = 32'b101001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [21] = 32'b101001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [22] = 32'b101001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [23] = 32'b101001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [24] = 32'b101001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [25] = 32'b101001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [26] = 32'b101001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [27] = 32'b101001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [28] = 32'b101001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [29] = 32'b101001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [30] = 32'b101001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r135 [31] = 32'b101001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [0] = 32'b101010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [1] = 32'b101010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [2] = 32'b101010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [3] = 32'b101010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [4] = 32'b101010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [5] = 32'b101010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [6] = 32'b101010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [7] = 32'b101010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [8] = 32'b101010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [9] = 32'b101010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [10] = 32'b101010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [11] = 32'b101010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [12] = 32'b101010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [13] = 32'b101010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [14] = 32'b101010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [15] = 32'b101010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [16] = 32'b101010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [17] = 32'b101010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [18] = 32'b101010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [19] = 32'b101010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [20] = 32'b101010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [21] = 32'b101010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [22] = 32'b101010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [23] = 32'b101010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [24] = 32'b101010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [25] = 32'b101010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [26] = 32'b101010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [27] = 32'b101010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [28] = 32'b101010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [29] = 32'b101010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [30] = 32'b101010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r134 [31] = 32'b101010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [0] = 32'b101010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [1] = 32'b101010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [2] = 32'b101010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [3] = 32'b101010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [4] = 32'b101010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [5] = 32'b101010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [6] = 32'b101010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [7] = 32'b101010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [8] = 32'b101010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [9] = 32'b101010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [10] = 32'b101010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [11] = 32'b101010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [12] = 32'b101010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [13] = 32'b101010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [14] = 32'b101010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [15] = 32'b101010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [16] = 32'b101010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [17] = 32'b101010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [18] = 32'b101010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [19] = 32'b101010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [20] = 32'b101010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [21] = 32'b101010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [22] = 32'b101010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [23] = 32'b101010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [24] = 32'b101010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [25] = 32'b101010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [26] = 32'b101010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [27] = 32'b101010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [28] = 32'b101010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [29] = 32'b101010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [30] = 32'b101010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r135 [31] = 32'b101010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [0] = 32'b101011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [1] = 32'b101011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [2] = 32'b101011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [3] = 32'b101011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [4] = 32'b101011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [5] = 32'b101011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [6] = 32'b101011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [7] = 32'b101011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [8] = 32'b101011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [9] = 32'b101011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [10] = 32'b101011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [11] = 32'b101011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [12] = 32'b101011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [13] = 32'b101011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [14] = 32'b101011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [15] = 32'b101011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [16] = 32'b101011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [17] = 32'b101011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [18] = 32'b101011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [19] = 32'b101011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [20] = 32'b101011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [21] = 32'b101011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [22] = 32'b101011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [23] = 32'b101011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [24] = 32'b101011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [25] = 32'b101011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [26] = 32'b101011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [27] = 32'b101011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [28] = 32'b101011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [29] = 32'b101011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [30] = 32'b101011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r134 [31] = 32'b101011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [0] = 32'b101011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [1] = 32'b101011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [2] = 32'b101011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [3] = 32'b101011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [4] = 32'b101011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [5] = 32'b101011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [6] = 32'b101011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [7] = 32'b101011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [8] = 32'b101011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [9] = 32'b101011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [10] = 32'b101011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [11] = 32'b101011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [12] = 32'b101011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [13] = 32'b101011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [14] = 32'b101011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [15] = 32'b101011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [16] = 32'b101011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [17] = 32'b101011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [18] = 32'b101011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [19] = 32'b101011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [20] = 32'b101011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [21] = 32'b101011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [22] = 32'b101011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [23] = 32'b101011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [24] = 32'b101011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [25] = 32'b101011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [26] = 32'b101011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [27] = 32'b101011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [28] = 32'b101011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [29] = 32'b101011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [30] = 32'b101011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r135 [31] = 32'b101011_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [0] = 32'b101100_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [1] = 32'b101100_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [2] = 32'b101100_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [3] = 32'b101100_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [4] = 32'b101100_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [5] = 32'b101100_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [6] = 32'b101100_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [7] = 32'b101100_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [8] = 32'b101100_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [9] = 32'b101100_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [10] = 32'b101100_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [11] = 32'b101100_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [12] = 32'b101100_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [13] = 32'b101100_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [14] = 32'b101100_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [15] = 32'b101100_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [16] = 32'b101100_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [17] = 32'b101100_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [18] = 32'b101100_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [19] = 32'b101100_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [20] = 32'b101100_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [21] = 32'b101100_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [22] = 32'b101100_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [23] = 32'b101100_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [24] = 32'b101100_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [25] = 32'b101100_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [26] = 32'b101100_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [27] = 32'b101100_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [28] = 32'b101100_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [29] = 32'b101100_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [30] = 32'b101100_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r134 [31] = 32'b101100_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [0] = 32'b101100_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [1] = 32'b101100_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [2] = 32'b101100_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [3] = 32'b101100_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [4] = 32'b101100_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [5] = 32'b101100_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [6] = 32'b101100_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [7] = 32'b101100_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [8] = 32'b101100_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [9] = 32'b101100_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [10] = 32'b101100_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [11] = 32'b101100_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [12] = 32'b101100_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [13] = 32'b101100_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [14] = 32'b101100_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [15] = 32'b101100_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [16] = 32'b101100_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [17] = 32'b101100_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [18] = 32'b101100_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [19] = 32'b101100_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [20] = 32'b101100_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [21] = 32'b101100_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [22] = 32'b101100_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [23] = 32'b101100_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [24] = 32'b101100_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [25] = 32'b101100_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [26] = 32'b101100_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [27] = 32'b101100_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [28] = 32'b101100_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [29] = 32'b101100_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [30] = 32'b101100_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r135 [31] = 32'b101100_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [0] = 32'b101101_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [1] = 32'b101101_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [2] = 32'b101101_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [3] = 32'b101101_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [4] = 32'b101101_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [5] = 32'b101101_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [6] = 32'b101101_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [7] = 32'b101101_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [8] = 32'b101101_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [9] = 32'b101101_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [10] = 32'b101101_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [11] = 32'b101101_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [12] = 32'b101101_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [13] = 32'b101101_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [14] = 32'b101101_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [15] = 32'b101101_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [16] = 32'b101101_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [17] = 32'b101101_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [18] = 32'b101101_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [19] = 32'b101101_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [20] = 32'b101101_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [21] = 32'b101101_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [22] = 32'b101101_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [23] = 32'b101101_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [24] = 32'b101101_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [25] = 32'b101101_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [26] = 32'b101101_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [27] = 32'b101101_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [28] = 32'b101101_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [29] = 32'b101101_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [30] = 32'b101101_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r134 [31] = 32'b101101_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [0] = 32'b101101_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [1] = 32'b101101_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [2] = 32'b101101_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [3] = 32'b101101_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [4] = 32'b101101_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [5] = 32'b101101_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [6] = 32'b101101_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [7] = 32'b101101_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [8] = 32'b101101_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [9] = 32'b101101_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [10] = 32'b101101_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [11] = 32'b101101_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [12] = 32'b101101_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [13] = 32'b101101_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [14] = 32'b101101_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [15] = 32'b101101_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [16] = 32'b101101_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [17] = 32'b101101_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [18] = 32'b101101_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [19] = 32'b101101_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [20] = 32'b101101_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [21] = 32'b101101_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [22] = 32'b101101_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [23] = 32'b101101_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [24] = 32'b101101_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [25] = 32'b101101_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [26] = 32'b101101_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [27] = 32'b101101_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [28] = 32'b101101_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [29] = 32'b101101_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [30] = 32'b101101_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r135 [31] = 32'b101101_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [0] = 32'b101110_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [1] = 32'b101110_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [2] = 32'b101110_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [3] = 32'b101110_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [4] = 32'b101110_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [5] = 32'b101110_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [6] = 32'b101110_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [7] = 32'b101110_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [8] = 32'b101110_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [9] = 32'b101110_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [10] = 32'b101110_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [11] = 32'b101110_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [12] = 32'b101110_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [13] = 32'b101110_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [14] = 32'b101110_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [15] = 32'b101110_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [16] = 32'b101110_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [17] = 32'b101110_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [18] = 32'b101110_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [19] = 32'b101110_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [20] = 32'b101110_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [21] = 32'b101110_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [22] = 32'b101110_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [23] = 32'b101110_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [24] = 32'b101110_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [25] = 32'b101110_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [26] = 32'b101110_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [27] = 32'b101110_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [28] = 32'b101110_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [29] = 32'b101110_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [30] = 32'b101110_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r134 [31] = 32'b101110_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [0] = 32'b101110_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [1] = 32'b101110_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [2] = 32'b101110_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [3] = 32'b101110_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [4] = 32'b101110_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [5] = 32'b101110_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [6] = 32'b101110_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [7] = 32'b101110_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [8] = 32'b101110_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [9] = 32'b101110_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [10] = 32'b101110_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [11] = 32'b101110_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [12] = 32'b101110_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [13] = 32'b101110_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [14] = 32'b101110_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [15] = 32'b101110_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [16] = 32'b101110_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [17] = 32'b101110_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [18] = 32'b101110_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [19] = 32'b101110_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [20] = 32'b101110_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [21] = 32'b101110_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [22] = 32'b101110_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [23] = 32'b101110_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [24] = 32'b101110_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [25] = 32'b101110_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [26] = 32'b101110_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [27] = 32'b101110_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [28] = 32'b101110_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [29] = 32'b101110_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [30] = 32'b101110_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r135 [31] = 32'b101110_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [0] = 32'b101111_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [1] = 32'b101111_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [2] = 32'b101111_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [3] = 32'b101111_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [4] = 32'b101111_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [5] = 32'b101111_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [6] = 32'b101111_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [7] = 32'b101111_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [8] = 32'b101111_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [9] = 32'b101111_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [10] = 32'b101111_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [11] = 32'b101111_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [12] = 32'b101111_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [13] = 32'b101111_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [14] = 32'b101111_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [15] = 32'b101111_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [16] = 32'b101111_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [17] = 32'b101111_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [18] = 32'b101111_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [19] = 32'b101111_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [20] = 32'b101111_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [21] = 32'b101111_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [22] = 32'b101111_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [23] = 32'b101111_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [24] = 32'b101111_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [25] = 32'b101111_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [26] = 32'b101111_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [27] = 32'b101111_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [28] = 32'b101111_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [29] = 32'b101111_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [30] = 32'b101111_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r134 [31] = 32'b101111_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [0] = 32'b101111_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [1] = 32'b101111_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [2] = 32'b101111_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [3] = 32'b101111_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [4] = 32'b101111_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [5] = 32'b101111_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [6] = 32'b101111_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [7] = 32'b101111_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [8] = 32'b101111_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [9] = 32'b101111_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [10] = 32'b101111_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [11] = 32'b101111_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [12] = 32'b101111_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [13] = 32'b101111_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [14] = 32'b101111_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [15] = 32'b101111_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [16] = 32'b101111_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [17] = 32'b101111_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [18] = 32'b101111_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [19] = 32'b101111_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [20] = 32'b101111_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [21] = 32'b101111_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [22] = 32'b101111_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [23] = 32'b101111_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [24] = 32'b101111_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [25] = 32'b101111_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [26] = 32'b101111_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [27] = 32'b101111_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [28] = 32'b101111_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [29] = 32'b101111_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [30] = 32'b101111_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r135 [31] = 32'b101111_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [0] = 32'b110000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [1] = 32'b110000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [2] = 32'b110000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [3] = 32'b110000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [4] = 32'b110000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [5] = 32'b110000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [6] = 32'b110000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [7] = 32'b110000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [8] = 32'b110000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [9] = 32'b110000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [10] = 32'b110000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [11] = 32'b110000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [12] = 32'b110000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [13] = 32'b110000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [14] = 32'b110000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [15] = 32'b110000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [16] = 32'b110000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [17] = 32'b110000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [18] = 32'b110000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [19] = 32'b110000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [20] = 32'b110000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [21] = 32'b110000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [22] = 32'b110000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [23] = 32'b110000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [24] = 32'b110000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [25] = 32'b110000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [26] = 32'b110000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [27] = 32'b110000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [28] = 32'b110000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [29] = 32'b110000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [30] = 32'b110000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r134 [31] = 32'b110000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [0] = 32'b110000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [1] = 32'b110000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [2] = 32'b110000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [3] = 32'b110000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [4] = 32'b110000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [5] = 32'b110000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [6] = 32'b110000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [7] = 32'b110000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [8] = 32'b110000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [9] = 32'b110000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [10] = 32'b110000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [11] = 32'b110000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [12] = 32'b110000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [13] = 32'b110000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [14] = 32'b110000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [15] = 32'b110000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [16] = 32'b110000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [17] = 32'b110000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [18] = 32'b110000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [19] = 32'b110000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [20] = 32'b110000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [21] = 32'b110000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [22] = 32'b110000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [23] = 32'b110000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [24] = 32'b110000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [25] = 32'b110000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [26] = 32'b110000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [27] = 32'b110000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [28] = 32'b110000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [29] = 32'b110000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [30] = 32'b110000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r135 [31] = 32'b110000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [0] = 32'b110001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [1] = 32'b110001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [2] = 32'b110001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [3] = 32'b110001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [4] = 32'b110001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [5] = 32'b110001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [6] = 32'b110001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [7] = 32'b110001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [8] = 32'b110001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [9] = 32'b110001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [10] = 32'b110001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [11] = 32'b110001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [12] = 32'b110001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [13] = 32'b110001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [14] = 32'b110001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [15] = 32'b110001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [16] = 32'b110001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [17] = 32'b110001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [18] = 32'b110001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [19] = 32'b110001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [20] = 32'b110001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [21] = 32'b110001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [22] = 32'b110001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [23] = 32'b110001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [24] = 32'b110001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [25] = 32'b110001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [26] = 32'b110001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [27] = 32'b110001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [28] = 32'b110001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [29] = 32'b110001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [30] = 32'b110001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r134 [31] = 32'b110001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [0] = 32'b110001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [1] = 32'b110001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [2] = 32'b110001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [3] = 32'b110001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [4] = 32'b110001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [5] = 32'b110001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [6] = 32'b110001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [7] = 32'b110001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [8] = 32'b110001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [9] = 32'b110001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [10] = 32'b110001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [11] = 32'b110001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [12] = 32'b110001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [13] = 32'b110001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [14] = 32'b110001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [15] = 32'b110001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [16] = 32'b110001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [17] = 32'b110001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [18] = 32'b110001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [19] = 32'b110001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [20] = 32'b110001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [21] = 32'b110001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [22] = 32'b110001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [23] = 32'b110001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [24] = 32'b110001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [25] = 32'b110001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [26] = 32'b110001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [27] = 32'b110001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [28] = 32'b110001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [29] = 32'b110001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [30] = 32'b110001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r135 [31] = 32'b110001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [0] = 32'b110010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [1] = 32'b110010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [2] = 32'b110010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [3] = 32'b110010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [4] = 32'b110010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [5] = 32'b110010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [6] = 32'b110010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [7] = 32'b110010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [8] = 32'b110010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [9] = 32'b110010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [10] = 32'b110010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [11] = 32'b110010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [12] = 32'b110010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [13] = 32'b110010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [14] = 32'b110010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [15] = 32'b110010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [16] = 32'b110010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [17] = 32'b110010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [18] = 32'b110010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [19] = 32'b110010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [20] = 32'b110010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [21] = 32'b110010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [22] = 32'b110010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [23] = 32'b110010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [24] = 32'b110010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [25] = 32'b110010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [26] = 32'b110010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [27] = 32'b110010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [28] = 32'b110010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [29] = 32'b110010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [30] = 32'b110010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r134 [31] = 32'b110010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [0] = 32'b110010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [1] = 32'b110010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [2] = 32'b110010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [3] = 32'b110010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [4] = 32'b110010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [5] = 32'b110010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [6] = 32'b110010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [7] = 32'b110010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [8] = 32'b110010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [9] = 32'b110010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [10] = 32'b110010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [11] = 32'b110010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [12] = 32'b110010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [13] = 32'b110010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [14] = 32'b110010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [15] = 32'b110010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [16] = 32'b110010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [17] = 32'b110010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [18] = 32'b110010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [19] = 32'b110010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [20] = 32'b110010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [21] = 32'b110010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [22] = 32'b110010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [23] = 32'b110010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [24] = 32'b110010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [25] = 32'b110010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [26] = 32'b110010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [27] = 32'b110010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [28] = 32'b110010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [29] = 32'b110010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [30] = 32'b110010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r135 [31] = 32'b110010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [0] = 32'b110011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [1] = 32'b110011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [2] = 32'b110011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [3] = 32'b110011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [4] = 32'b110011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [5] = 32'b110011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [6] = 32'b110011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [7] = 32'b110011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [8] = 32'b110011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [9] = 32'b110011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [10] = 32'b110011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [11] = 32'b110011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [12] = 32'b110011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [13] = 32'b110011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [14] = 32'b110011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [15] = 32'b110011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [16] = 32'b110011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [17] = 32'b110011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [18] = 32'b110011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [19] = 32'b110011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [20] = 32'b110011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [21] = 32'b110011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [22] = 32'b110011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [23] = 32'b110011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [24] = 32'b110011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [25] = 32'b110011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [26] = 32'b110011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [27] = 32'b110011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [28] = 32'b110011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [29] = 32'b110011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [30] = 32'b110011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r134 [31] = 32'b110011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [0] = 32'b110011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [1] = 32'b110011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [2] = 32'b110011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [3] = 32'b110011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [4] = 32'b110011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [5] = 32'b110011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [6] = 32'b110011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [7] = 32'b110011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [8] = 32'b110011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [9] = 32'b110011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [10] = 32'b110011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [11] = 32'b110011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [12] = 32'b110011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [13] = 32'b110011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [14] = 32'b110011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [15] = 32'b110011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [16] = 32'b110011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [17] = 32'b110011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [18] = 32'b110011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [19] = 32'b110011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [20] = 32'b110011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [21] = 32'b110011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [22] = 32'b110011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [23] = 32'b110011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [24] = 32'b110011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [25] = 32'b110011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [26] = 32'b110011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [27] = 32'b110011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [28] = 32'b110011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [29] = 32'b110011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [30] = 32'b110011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r135 [31] = 32'b110011_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [0] = 32'b110100_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [1] = 32'b110100_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [2] = 32'b110100_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [3] = 32'b110100_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [4] = 32'b110100_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [5] = 32'b110100_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [6] = 32'b110100_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [7] = 32'b110100_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [8] = 32'b110100_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [9] = 32'b110100_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [10] = 32'b110100_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [11] = 32'b110100_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [12] = 32'b110100_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [13] = 32'b110100_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [14] = 32'b110100_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [15] = 32'b110100_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [16] = 32'b110100_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [17] = 32'b110100_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [18] = 32'b110100_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [19] = 32'b110100_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [20] = 32'b110100_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [21] = 32'b110100_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [22] = 32'b110100_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [23] = 32'b110100_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [24] = 32'b110100_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [25] = 32'b110100_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [26] = 32'b110100_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [27] = 32'b110100_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [28] = 32'b110100_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [29] = 32'b110100_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [30] = 32'b110100_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r134 [31] = 32'b110100_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [0] = 32'b110100_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [1] = 32'b110100_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [2] = 32'b110100_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [3] = 32'b110100_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [4] = 32'b110100_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [5] = 32'b110100_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [6] = 32'b110100_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [7] = 32'b110100_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [8] = 32'b110100_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [9] = 32'b110100_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [10] = 32'b110100_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [11] = 32'b110100_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [12] = 32'b110100_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [13] = 32'b110100_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [14] = 32'b110100_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [15] = 32'b110100_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [16] = 32'b110100_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [17] = 32'b110100_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [18] = 32'b110100_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [19] = 32'b110100_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [20] = 32'b110100_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [21] = 32'b110100_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [22] = 32'b110100_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [23] = 32'b110100_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [24] = 32'b110100_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [25] = 32'b110100_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [26] = 32'b110100_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [27] = 32'b110100_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [28] = 32'b110100_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [29] = 32'b110100_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [30] = 32'b110100_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r135 [31] = 32'b110100_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [0] = 32'b110101_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [1] = 32'b110101_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [2] = 32'b110101_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [3] = 32'b110101_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [4] = 32'b110101_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [5] = 32'b110101_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [6] = 32'b110101_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [7] = 32'b110101_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [8] = 32'b110101_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [9] = 32'b110101_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [10] = 32'b110101_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [11] = 32'b110101_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [12] = 32'b110101_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [13] = 32'b110101_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [14] = 32'b110101_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [15] = 32'b110101_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [16] = 32'b110101_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [17] = 32'b110101_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [18] = 32'b110101_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [19] = 32'b110101_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [20] = 32'b110101_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [21] = 32'b110101_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [22] = 32'b110101_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [23] = 32'b110101_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [24] = 32'b110101_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [25] = 32'b110101_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [26] = 32'b110101_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [27] = 32'b110101_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [28] = 32'b110101_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [29] = 32'b110101_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [30] = 32'b110101_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r134 [31] = 32'b110101_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [0] = 32'b110101_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [1] = 32'b110101_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [2] = 32'b110101_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [3] = 32'b110101_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [4] = 32'b110101_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [5] = 32'b110101_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [6] = 32'b110101_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [7] = 32'b110101_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [8] = 32'b110101_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [9] = 32'b110101_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [10] = 32'b110101_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [11] = 32'b110101_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [12] = 32'b110101_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [13] = 32'b110101_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [14] = 32'b110101_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [15] = 32'b110101_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [16] = 32'b110101_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [17] = 32'b110101_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [18] = 32'b110101_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [19] = 32'b110101_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [20] = 32'b110101_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [21] = 32'b110101_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [22] = 32'b110101_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [23] = 32'b110101_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [24] = 32'b110101_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [25] = 32'b110101_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [26] = 32'b110101_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [27] = 32'b110101_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [28] = 32'b110101_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [29] = 32'b110101_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [30] = 32'b110101_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r135 [31] = 32'b110101_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [0] = 32'b110110_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [1] = 32'b110110_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [2] = 32'b110110_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [3] = 32'b110110_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [4] = 32'b110110_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [5] = 32'b110110_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [6] = 32'b110110_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [7] = 32'b110110_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [8] = 32'b110110_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [9] = 32'b110110_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [10] = 32'b110110_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [11] = 32'b110110_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [12] = 32'b110110_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [13] = 32'b110110_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [14] = 32'b110110_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [15] = 32'b110110_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [16] = 32'b110110_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [17] = 32'b110110_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [18] = 32'b110110_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [19] = 32'b110110_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [20] = 32'b110110_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [21] = 32'b110110_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [22] = 32'b110110_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [23] = 32'b110110_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [24] = 32'b110110_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [25] = 32'b110110_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [26] = 32'b110110_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [27] = 32'b110110_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [28] = 32'b110110_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [29] = 32'b110110_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [30] = 32'b110110_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r134 [31] = 32'b110110_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [0] = 32'b110110_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [1] = 32'b110110_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [2] = 32'b110110_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [3] = 32'b110110_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [4] = 32'b110110_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [5] = 32'b110110_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [6] = 32'b110110_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [7] = 32'b110110_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [8] = 32'b110110_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [9] = 32'b110110_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [10] = 32'b110110_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [11] = 32'b110110_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [12] = 32'b110110_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [13] = 32'b110110_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [14] = 32'b110110_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [15] = 32'b110110_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [16] = 32'b110110_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [17] = 32'b110110_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [18] = 32'b110110_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [19] = 32'b110110_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [20] = 32'b110110_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [21] = 32'b110110_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [22] = 32'b110110_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [23] = 32'b110110_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [24] = 32'b110110_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [25] = 32'b110110_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [26] = 32'b110110_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [27] = 32'b110110_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [28] = 32'b110110_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [29] = 32'b110110_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [30] = 32'b110110_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r135 [31] = 32'b110110_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [0] = 32'b110111_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [1] = 32'b110111_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [2] = 32'b110111_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [3] = 32'b110111_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [4] = 32'b110111_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [5] = 32'b110111_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [6] = 32'b110111_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [7] = 32'b110111_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [8] = 32'b110111_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [9] = 32'b110111_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [10] = 32'b110111_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [11] = 32'b110111_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [12] = 32'b110111_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [13] = 32'b110111_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [14] = 32'b110111_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [15] = 32'b110111_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [16] = 32'b110111_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [17] = 32'b110111_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [18] = 32'b110111_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [19] = 32'b110111_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [20] = 32'b110111_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [21] = 32'b110111_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [22] = 32'b110111_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [23] = 32'b110111_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [24] = 32'b110111_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [25] = 32'b110111_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [26] = 32'b110111_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [27] = 32'b110111_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [28] = 32'b110111_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [29] = 32'b110111_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [30] = 32'b110111_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r134 [31] = 32'b110111_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [0] = 32'b110111_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [1] = 32'b110111_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [2] = 32'b110111_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [3] = 32'b110111_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [4] = 32'b110111_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [5] = 32'b110111_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [6] = 32'b110111_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [7] = 32'b110111_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [8] = 32'b110111_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [9] = 32'b110111_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [10] = 32'b110111_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [11] = 32'b110111_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [12] = 32'b110111_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [13] = 32'b110111_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [14] = 32'b110111_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [15] = 32'b110111_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [16] = 32'b110111_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [17] = 32'b110111_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [18] = 32'b110111_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [19] = 32'b110111_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [20] = 32'b110111_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [21] = 32'b110111_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [22] = 32'b110111_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [23] = 32'b110111_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [24] = 32'b110111_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [25] = 32'b110111_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [26] = 32'b110111_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [27] = 32'b110111_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [28] = 32'b110111_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [29] = 32'b110111_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [30] = 32'b110111_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r135 [31] = 32'b110111_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [0] = 32'b111000_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [1] = 32'b111000_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [2] = 32'b111000_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [3] = 32'b111000_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [4] = 32'b111000_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [5] = 32'b111000_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [6] = 32'b111000_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [7] = 32'b111000_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [8] = 32'b111000_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [9] = 32'b111000_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [10] = 32'b111000_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [11] = 32'b111000_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [12] = 32'b111000_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [13] = 32'b111000_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [14] = 32'b111000_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [15] = 32'b111000_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [16] = 32'b111000_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [17] = 32'b111000_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [18] = 32'b111000_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [19] = 32'b111000_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [20] = 32'b111000_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [21] = 32'b111000_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [22] = 32'b111000_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [23] = 32'b111000_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [24] = 32'b111000_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [25] = 32'b111000_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [26] = 32'b111000_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [27] = 32'b111000_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [28] = 32'b111000_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [29] = 32'b111000_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [30] = 32'b111000_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r134 [31] = 32'b111000_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [0] = 32'b111000_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [1] = 32'b111000_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [2] = 32'b111000_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [3] = 32'b111000_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [4] = 32'b111000_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [5] = 32'b111000_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [6] = 32'b111000_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [7] = 32'b111000_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [8] = 32'b111000_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [9] = 32'b111000_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [10] = 32'b111000_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [11] = 32'b111000_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [12] = 32'b111000_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [13] = 32'b111000_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [14] = 32'b111000_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [15] = 32'b111000_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [16] = 32'b111000_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [17] = 32'b111000_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [18] = 32'b111000_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [19] = 32'b111000_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [20] = 32'b111000_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [21] = 32'b111000_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [22] = 32'b111000_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [23] = 32'b111000_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [24] = 32'b111000_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [25] = 32'b111000_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [26] = 32'b111000_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [27] = 32'b111000_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [28] = 32'b111000_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [29] = 32'b111000_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [30] = 32'b111000_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r135 [31] = 32'b111000_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [0] = 32'b111001_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [1] = 32'b111001_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [2] = 32'b111001_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [3] = 32'b111001_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [4] = 32'b111001_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [5] = 32'b111001_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [6] = 32'b111001_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [7] = 32'b111001_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [8] = 32'b111001_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [9] = 32'b111001_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [10] = 32'b111001_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [11] = 32'b111001_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [12] = 32'b111001_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [13] = 32'b111001_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [14] = 32'b111001_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [15] = 32'b111001_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [16] = 32'b111001_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [17] = 32'b111001_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [18] = 32'b111001_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [19] = 32'b111001_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [20] = 32'b111001_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [21] = 32'b111001_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [22] = 32'b111001_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [23] = 32'b111001_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [24] = 32'b111001_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [25] = 32'b111001_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [26] = 32'b111001_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [27] = 32'b111001_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [28] = 32'b111001_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [29] = 32'b111001_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [30] = 32'b111001_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r134 [31] = 32'b111001_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [0] = 32'b111001_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [1] = 32'b111001_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [2] = 32'b111001_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [3] = 32'b111001_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [4] = 32'b111001_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [5] = 32'b111001_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [6] = 32'b111001_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [7] = 32'b111001_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [8] = 32'b111001_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [9] = 32'b111001_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [10] = 32'b111001_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [11] = 32'b111001_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [12] = 32'b111001_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [13] = 32'b111001_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [14] = 32'b111001_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [15] = 32'b111001_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [16] = 32'b111001_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [17] = 32'b111001_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [18] = 32'b111001_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [19] = 32'b111001_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [20] = 32'b111001_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [21] = 32'b111001_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [22] = 32'b111001_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [23] = 32'b111001_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [24] = 32'b111001_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [25] = 32'b111001_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [26] = 32'b111001_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [27] = 32'b111001_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [28] = 32'b111001_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [29] = 32'b111001_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [30] = 32'b111001_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r135 [31] = 32'b111001_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [0] = 32'b111010_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [1] = 32'b111010_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [2] = 32'b111010_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [3] = 32'b111010_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [4] = 32'b111010_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [5] = 32'b111010_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [6] = 32'b111010_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [7] = 32'b111010_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [8] = 32'b111010_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [9] = 32'b111010_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [10] = 32'b111010_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [11] = 32'b111010_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [12] = 32'b111010_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [13] = 32'b111010_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [14] = 32'b111010_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [15] = 32'b111010_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [16] = 32'b111010_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [17] = 32'b111010_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [18] = 32'b111010_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [19] = 32'b111010_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [20] = 32'b111010_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [21] = 32'b111010_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [22] = 32'b111010_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [23] = 32'b111010_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [24] = 32'b111010_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [25] = 32'b111010_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [26] = 32'b111010_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [27] = 32'b111010_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [28] = 32'b111010_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [29] = 32'b111010_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [30] = 32'b111010_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r134 [31] = 32'b111010_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [0] = 32'b111010_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [1] = 32'b111010_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [2] = 32'b111010_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [3] = 32'b111010_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [4] = 32'b111010_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [5] = 32'b111010_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [6] = 32'b111010_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [7] = 32'b111010_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [8] = 32'b111010_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [9] = 32'b111010_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [10] = 32'b111010_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [11] = 32'b111010_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [12] = 32'b111010_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [13] = 32'b111010_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [14] = 32'b111010_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [15] = 32'b111010_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [16] = 32'b111010_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [17] = 32'b111010_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [18] = 32'b111010_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [19] = 32'b111010_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [20] = 32'b111010_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [21] = 32'b111010_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [22] = 32'b111010_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [23] = 32'b111010_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [24] = 32'b111010_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [25] = 32'b111010_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [26] = 32'b111010_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [27] = 32'b111010_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [28] = 32'b111010_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [29] = 32'b111010_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [30] = 32'b111010_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r135 [31] = 32'b111010_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [0] = 32'b111011_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [1] = 32'b111011_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [2] = 32'b111011_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [3] = 32'b111011_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [4] = 32'b111011_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [5] = 32'b111011_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [6] = 32'b111011_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [7] = 32'b111011_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [8] = 32'b111011_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [9] = 32'b111011_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [10] = 32'b111011_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [11] = 32'b111011_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [12] = 32'b111011_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [13] = 32'b111011_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [14] = 32'b111011_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [15] = 32'b111011_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [16] = 32'b111011_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [17] = 32'b111011_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [18] = 32'b111011_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [19] = 32'b111011_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [20] = 32'b111011_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [21] = 32'b111011_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [22] = 32'b111011_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [23] = 32'b111011_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [24] = 32'b111011_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [25] = 32'b111011_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [26] = 32'b111011_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [27] = 32'b111011_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [28] = 32'b111011_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [29] = 32'b111011_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [30] = 32'b111011_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r134 [31] = 32'b111011_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [0] = 32'b111011_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [1] = 32'b111011_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [2] = 32'b111011_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [3] = 32'b111011_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [4] = 32'b111011_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [5] = 32'b111011_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [6] = 32'b111011_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [7] = 32'b111011_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [8] = 32'b111011_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [9] = 32'b111011_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [10] = 32'b111011_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [11] = 32'b111011_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [12] = 32'b111011_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [13] = 32'b111011_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [14] = 32'b111011_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [15] = 32'b111011_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [16] = 32'b111011_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [17] = 32'b111011_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [18] = 32'b111011_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [19] = 32'b111011_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [20] = 32'b111011_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [21] = 32'b111011_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [22] = 32'b111011_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [23] = 32'b111011_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [24] = 32'b111011_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [25] = 32'b111011_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [26] = 32'b111011_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [27] = 32'b111011_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [28] = 32'b111011_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [29] = 32'b111011_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [30] = 32'b111011_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r135 [31] = 32'b111011_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [0] = 32'b111100_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [1] = 32'b111100_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [2] = 32'b111100_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [3] = 32'b111100_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [4] = 32'b111100_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [5] = 32'b111100_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [6] = 32'b111100_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [7] = 32'b111100_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [8] = 32'b111100_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [9] = 32'b111100_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [10] = 32'b111100_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [11] = 32'b111100_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [12] = 32'b111100_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [13] = 32'b111100_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [14] = 32'b111100_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [15] = 32'b111100_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [16] = 32'b111100_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [17] = 32'b111100_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [18] = 32'b111100_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [19] = 32'b111100_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [20] = 32'b111100_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [21] = 32'b111100_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [22] = 32'b111100_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [23] = 32'b111100_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [24] = 32'b111100_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [25] = 32'b111100_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [26] = 32'b111100_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [27] = 32'b111100_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [28] = 32'b111100_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [29] = 32'b111100_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [30] = 32'b111100_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r134 [31] = 32'b111100_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [0] = 32'b111100_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [1] = 32'b111100_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [2] = 32'b111100_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [3] = 32'b111100_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [4] = 32'b111100_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [5] = 32'b111100_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [6] = 32'b111100_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [7] = 32'b111100_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [8] = 32'b111100_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [9] = 32'b111100_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [10] = 32'b111100_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [11] = 32'b111100_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [12] = 32'b111100_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [13] = 32'b111100_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [14] = 32'b111100_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [15] = 32'b111100_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [16] = 32'b111100_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [17] = 32'b111100_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [18] = 32'b111100_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [19] = 32'b111100_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [20] = 32'b111100_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [21] = 32'b111100_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [22] = 32'b111100_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [23] = 32'b111100_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [24] = 32'b111100_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [25] = 32'b111100_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [26] = 32'b111100_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [27] = 32'b111100_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [28] = 32'b111100_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [29] = 32'b111100_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [30] = 32'b111100_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r135 [31] = 32'b111100_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [0] = 32'b111101_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [1] = 32'b111101_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [2] = 32'b111101_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [3] = 32'b111101_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [4] = 32'b111101_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [5] = 32'b111101_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [6] = 32'b111101_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [7] = 32'b111101_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [8] = 32'b111101_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [9] = 32'b111101_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [10] = 32'b111101_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [11] = 32'b111101_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [12] = 32'b111101_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [13] = 32'b111101_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [14] = 32'b111101_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [15] = 32'b111101_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [16] = 32'b111101_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [17] = 32'b111101_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [18] = 32'b111101_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [19] = 32'b111101_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [20] = 32'b111101_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [21] = 32'b111101_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [22] = 32'b111101_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [23] = 32'b111101_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [24] = 32'b111101_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [25] = 32'b111101_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [26] = 32'b111101_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [27] = 32'b111101_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [28] = 32'b111101_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [29] = 32'b111101_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [30] = 32'b111101_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r134 [31] = 32'b111101_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [0] = 32'b111101_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [1] = 32'b111101_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [2] = 32'b111101_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [3] = 32'b111101_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [4] = 32'b111101_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [5] = 32'b111101_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [6] = 32'b111101_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [7] = 32'b111101_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [8] = 32'b111101_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [9] = 32'b111101_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [10] = 32'b111101_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [11] = 32'b111101_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [12] = 32'b111101_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [13] = 32'b111101_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [14] = 32'b111101_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [15] = 32'b111101_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [16] = 32'b111101_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [17] = 32'b111101_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [18] = 32'b111101_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [19] = 32'b111101_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [20] = 32'b111101_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [21] = 32'b111101_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [22] = 32'b111101_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [23] = 32'b111101_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [24] = 32'b111101_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [25] = 32'b111101_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [26] = 32'b111101_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [27] = 32'b111101_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [28] = 32'b111101_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [29] = 32'b111101_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [30] = 32'b111101_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r135 [31] = 32'b111101_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [0] = 32'b111110_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [1] = 32'b111110_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [2] = 32'b111110_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [3] = 32'b111110_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [4] = 32'b111110_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [5] = 32'b111110_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [6] = 32'b111110_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [7] = 32'b111110_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [8] = 32'b111110_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [9] = 32'b111110_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [10] = 32'b111110_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [11] = 32'b111110_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [12] = 32'b111110_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [13] = 32'b111110_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [14] = 32'b111110_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [15] = 32'b111110_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [16] = 32'b111110_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [17] = 32'b111110_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [18] = 32'b111110_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [19] = 32'b111110_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [20] = 32'b111110_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [21] = 32'b111110_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [22] = 32'b111110_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [23] = 32'b111110_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [24] = 32'b111110_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [25] = 32'b111110_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [26] = 32'b111110_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [27] = 32'b111110_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [28] = 32'b111110_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [29] = 32'b111110_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [30] = 32'b111110_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r134 [31] = 32'b111110_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [0] = 32'b111110_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [1] = 32'b111110_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [2] = 32'b111110_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [3] = 32'b111110_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [4] = 32'b111110_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [5] = 32'b111110_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [6] = 32'b111110_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [7] = 32'b111110_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [8] = 32'b111110_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [9] = 32'b111110_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [10] = 32'b111110_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [11] = 32'b111110_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [12] = 32'b111110_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [13] = 32'b111110_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [14] = 32'b111110_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [15] = 32'b111110_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [16] = 32'b111110_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [17] = 32'b111110_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [18] = 32'b111110_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [19] = 32'b111110_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [20] = 32'b111110_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [21] = 32'b111110_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [22] = 32'b111110_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [23] = 32'b111110_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [24] = 32'b111110_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [25] = 32'b111110_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [26] = 32'b111110_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [27] = 32'b111110_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [28] = 32'b111110_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [29] = 32'b111110_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [30] = 32'b111110_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r135 [31] = 32'b111110_11111__0_1000_0000_0000;
            // Stream 0 Destination address
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [0] = 32'b111111_00000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [1] = 32'b111111_00001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [2] = 32'b111111_00010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [3] = 32'b111111_00011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [4] = 32'b111111_00100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [5] = 32'b111111_00101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [6] = 32'b111111_00110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [7] = 32'b111111_00111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [8] = 32'b111111_01000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [9] = 32'b111111_01001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [10] = 32'b111111_01010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [11] = 32'b111111_01011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [12] = 32'b111111_01100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [13] = 32'b111111_01101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [14] = 32'b111111_01110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [15] = 32'b111111_01111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [16] = 32'b111111_10000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [17] = 32'b111111_10001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [18] = 32'b111111_10010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [19] = 32'b111111_10011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [20] = 32'b111111_10100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [21] = 32'b111111_10101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [22] = 32'b111111_10110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [23] = 32'b111111_10111__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [24] = 32'b111111_11000__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [25] = 32'b111111_11001__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [26] = 32'b111111_11010__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [27] = 32'b111111_11011__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [28] = 32'b111111_11100__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [29] = 32'b111111_11101__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [30] = 32'b111111_11110__0_0000_1000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r134 [31] = 32'b111111_11111__0_0000_1000_0000;
            // Stream 1 Destination address
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [0] = 32'b111111_00000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [1] = 32'b111111_00001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [2] = 32'b111111_00010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [3] = 32'b111111_00011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [4] = 32'b111111_00100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [5] = 32'b111111_00101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [6] = 32'b111111_00110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [7] = 32'b111111_00111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [8] = 32'b111111_01000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [9] = 32'b111111_01001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [10] = 32'b111111_01010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [11] = 32'b111111_01011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [12] = 32'b111111_01100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [13] = 32'b111111_01101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [14] = 32'b111111_01110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [15] = 32'b111111_01111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [16] = 32'b111111_10000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [17] = 32'b111111_10001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [18] = 32'b111111_10010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [19] = 32'b111111_10011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [20] = 32'b111111_10100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [21] = 32'b111111_10101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [22] = 32'b111111_10110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [23] = 32'b111111_10111__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [24] = 32'b111111_11000__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [25] = 32'b111111_11001__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [26] = 32'b111111_11010__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [27] = 32'b111111_11011__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [28] = 32'b111111_11100__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [29] = 32'b111111_11101__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [30] = 32'b111111_11110__0_1000_0000_0000;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r135 [31] = 32'b111111_11111__0_1000_0000_0000;

            // ##################################################
            // DMA Type and length of stream

            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r132 [31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__lane_r133 [31][15:0]  = numOfTypes;

            // ##################################################
            // Enable Stack bus streams


            // ##################################################
            // Enable and set transfer type

            repeat(10) @(negedge clk); 

            // Enable
            force pe_array_inst.pe_inst[0].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__rs0[0]           = 1'b1;

            // Operation
            force pe_array_inst.pe_inst[0].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[4].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[5].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[6].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[7].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[8].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[9].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[10].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[11].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[12].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[13].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[14].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[15].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[16].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[17].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[18].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[19].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[20].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[21].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[22].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[23].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[24].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[25].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[26].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[27].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[28].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[29].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[30].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[31].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[32].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[33].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[34].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[35].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[36].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[37].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[38].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[39].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[40].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[41].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[42].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[43].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[44].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[45].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[46].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[47].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[48].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[49].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[50].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[51].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[52].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[53].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[54].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[55].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[56].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[57].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[58].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[59].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[60].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[61].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[62].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;
            force pe_array_inst.pe_inst[63].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM ;

            repeat(50) @(negedge clk);