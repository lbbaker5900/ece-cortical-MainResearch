
  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[0].mgr__sys__allSynchronized   =  GenStackBus[0].sys__pe__allSynchronized                                ; 
  assign GenStackBus[0].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[0].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[0].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[0].sys__mgr__ready             ; 
  assign GenStackBus[0].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[0].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[1].mgr__sys__allSynchronized   =  GenStackBus[1].sys__pe__allSynchronized                                ; 
  assign GenStackBus[1].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[1].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[1].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[1].sys__mgr__ready             ; 
  assign GenStackBus[1].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[1].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[2].mgr__sys__allSynchronized   =  GenStackBus[2].sys__pe__allSynchronized                                ; 
  assign GenStackBus[2].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[2].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[2].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[2].sys__mgr__ready             ; 
  assign GenStackBus[2].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[2].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[3].mgr__sys__allSynchronized   =  GenStackBus[3].sys__pe__allSynchronized                                ; 
  assign GenStackBus[3].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[3].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[3].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[3].sys__mgr__ready             ; 
  assign GenStackBus[3].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[3].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[4].mgr__sys__allSynchronized   =  GenStackBus[4].sys__pe__allSynchronized                                ; 
  assign GenStackBus[4].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[4].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[4].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[4].sys__mgr__ready             ; 
  assign GenStackBus[4].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[4].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[5].mgr__sys__allSynchronized   =  GenStackBus[5].sys__pe__allSynchronized                                ; 
  assign GenStackBus[5].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[5].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[5].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[5].sys__mgr__ready             ; 
  assign GenStackBus[5].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[5].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[6].mgr__sys__allSynchronized   =  GenStackBus[6].sys__pe__allSynchronized                                ; 
  assign GenStackBus[6].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[6].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[6].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[6].sys__mgr__ready             ; 
  assign GenStackBus[6].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[6].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[7].mgr__sys__allSynchronized   =  GenStackBus[7].sys__pe__allSynchronized                                ; 
  assign GenStackBus[7].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[7].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[7].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[7].sys__mgr__ready             ; 
  assign GenStackBus[7].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[7].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[8].mgr__sys__allSynchronized   =  GenStackBus[8].sys__pe__allSynchronized                                ; 
  assign GenStackBus[8].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[8].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[8].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[8].sys__mgr__ready             ; 
  assign GenStackBus[8].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[8].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[9].mgr__sys__allSynchronized   =  GenStackBus[9].sys__pe__allSynchronized                                ; 
  assign GenStackBus[9].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[9].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[9].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[9].sys__mgr__ready             ; 
  assign GenStackBus[9].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[9].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[10].mgr__sys__allSynchronized   =  GenStackBus[10].sys__pe__allSynchronized                                ; 
  assign GenStackBus[10].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[10].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[10].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[10].sys__mgr__ready             ; 
  assign GenStackBus[10].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[10].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[11].mgr__sys__allSynchronized   =  GenStackBus[11].sys__pe__allSynchronized                                ; 
  assign GenStackBus[11].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[11].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[11].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[11].sys__mgr__ready             ; 
  assign GenStackBus[11].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[11].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[12].mgr__sys__allSynchronized   =  GenStackBus[12].sys__pe__allSynchronized                                ; 
  assign GenStackBus[12].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[12].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[12].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[12].sys__mgr__ready             ; 
  assign GenStackBus[12].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[12].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[13].mgr__sys__allSynchronized   =  GenStackBus[13].sys__pe__allSynchronized                                ; 
  assign GenStackBus[13].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[13].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[13].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[13].sys__mgr__ready             ; 
  assign GenStackBus[13].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[13].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[14].mgr__sys__allSynchronized   =  GenStackBus[14].sys__pe__allSynchronized                                ; 
  assign GenStackBus[14].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[14].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[14].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[14].sys__mgr__ready             ; 
  assign GenStackBus[14].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[14].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[15].mgr__sys__allSynchronized   =  GenStackBus[15].sys__pe__allSynchronized                                ; 
  assign GenStackBus[15].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[15].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[15].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[15].sys__mgr__ready             ; 
  assign GenStackBus[15].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[15].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[16].mgr__sys__allSynchronized   =  GenStackBus[16].sys__pe__allSynchronized                                ; 
  assign GenStackBus[16].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[16].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[16].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[16].sys__mgr__ready             ; 
  assign GenStackBus[16].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[16].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[17].mgr__sys__allSynchronized   =  GenStackBus[17].sys__pe__allSynchronized                                ; 
  assign GenStackBus[17].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[17].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[17].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[17].sys__mgr__ready             ; 
  assign GenStackBus[17].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[17].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[18].mgr__sys__allSynchronized   =  GenStackBus[18].sys__pe__allSynchronized                                ; 
  assign GenStackBus[18].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[18].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[18].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[18].sys__mgr__ready             ; 
  assign GenStackBus[18].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[18].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[19].mgr__sys__allSynchronized   =  GenStackBus[19].sys__pe__allSynchronized                                ; 
  assign GenStackBus[19].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[19].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[19].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[19].sys__mgr__ready             ; 
  assign GenStackBus[19].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[19].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[20].mgr__sys__allSynchronized   =  GenStackBus[20].sys__pe__allSynchronized                                ; 
  assign GenStackBus[20].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[20].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[20].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[20].sys__mgr__ready             ; 
  assign GenStackBus[20].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[20].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[21].mgr__sys__allSynchronized   =  GenStackBus[21].sys__pe__allSynchronized                                ; 
  assign GenStackBus[21].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[21].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[21].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[21].sys__mgr__ready             ; 
  assign GenStackBus[21].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[21].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[22].mgr__sys__allSynchronized   =  GenStackBus[22].sys__pe__allSynchronized                                ; 
  assign GenStackBus[22].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[22].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[22].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[22].sys__mgr__ready             ; 
  assign GenStackBus[22].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[22].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[23].mgr__sys__allSynchronized   =  GenStackBus[23].sys__pe__allSynchronized                                ; 
  assign GenStackBus[23].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[23].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[23].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[23].sys__mgr__ready             ; 
  assign GenStackBus[23].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[23].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[24].mgr__sys__allSynchronized   =  GenStackBus[24].sys__pe__allSynchronized                                ; 
  assign GenStackBus[24].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[24].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[24].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[24].sys__mgr__ready             ; 
  assign GenStackBus[24].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[24].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[25].mgr__sys__allSynchronized   =  GenStackBus[25].sys__pe__allSynchronized                                ; 
  assign GenStackBus[25].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[25].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[25].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[25].sys__mgr__ready             ; 
  assign GenStackBus[25].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[25].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[26].mgr__sys__allSynchronized   =  GenStackBus[26].sys__pe__allSynchronized                                ; 
  assign GenStackBus[26].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[26].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[26].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[26].sys__mgr__ready             ; 
  assign GenStackBus[26].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[26].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[27].mgr__sys__allSynchronized   =  GenStackBus[27].sys__pe__allSynchronized                                ; 
  assign GenStackBus[27].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[27].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[27].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[27].sys__mgr__ready             ; 
  assign GenStackBus[27].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[27].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[28].mgr__sys__allSynchronized   =  GenStackBus[28].sys__pe__allSynchronized                                ; 
  assign GenStackBus[28].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[28].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[28].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[28].sys__mgr__ready             ; 
  assign GenStackBus[28].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[28].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[29].mgr__sys__allSynchronized   =  GenStackBus[29].sys__pe__allSynchronized                                ; 
  assign GenStackBus[29].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[29].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[29].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[29].sys__mgr__ready             ; 
  assign GenStackBus[29].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[29].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[30].mgr__sys__allSynchronized   =  GenStackBus[30].sys__pe__allSynchronized                                ; 
  assign GenStackBus[30].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[30].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[30].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[30].sys__mgr__ready             ; 
  assign GenStackBus[30].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[30].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[31].mgr__sys__allSynchronized   =  GenStackBus[31].sys__pe__allSynchronized                                ; 
  assign GenStackBus[31].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[31].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[31].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[31].sys__mgr__ready             ; 
  assign GenStackBus[31].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[31].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[32].mgr__sys__allSynchronized   =  GenStackBus[32].sys__pe__allSynchronized                                ; 
  assign GenStackBus[32].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[32].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[32].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[32].sys__mgr__ready             ; 
  assign GenStackBus[32].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[32].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[33].mgr__sys__allSynchronized   =  GenStackBus[33].sys__pe__allSynchronized                                ; 
  assign GenStackBus[33].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[33].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[33].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[33].sys__mgr__ready             ; 
  assign GenStackBus[33].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[33].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[34].mgr__sys__allSynchronized   =  GenStackBus[34].sys__pe__allSynchronized                                ; 
  assign GenStackBus[34].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[34].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[34].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[34].sys__mgr__ready             ; 
  assign GenStackBus[34].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[34].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[35].mgr__sys__allSynchronized   =  GenStackBus[35].sys__pe__allSynchronized                                ; 
  assign GenStackBus[35].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[35].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[35].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[35].sys__mgr__ready             ; 
  assign GenStackBus[35].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[35].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[36].mgr__sys__allSynchronized   =  GenStackBus[36].sys__pe__allSynchronized                                ; 
  assign GenStackBus[36].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[36].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[36].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[36].sys__mgr__ready             ; 
  assign GenStackBus[36].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[36].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[37].mgr__sys__allSynchronized   =  GenStackBus[37].sys__pe__allSynchronized                                ; 
  assign GenStackBus[37].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[37].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[37].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[37].sys__mgr__ready             ; 
  assign GenStackBus[37].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[37].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[38].mgr__sys__allSynchronized   =  GenStackBus[38].sys__pe__allSynchronized                                ; 
  assign GenStackBus[38].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[38].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[38].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[38].sys__mgr__ready             ; 
  assign GenStackBus[38].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[38].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[39].mgr__sys__allSynchronized   =  GenStackBus[39].sys__pe__allSynchronized                                ; 
  assign GenStackBus[39].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[39].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[39].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[39].sys__mgr__ready             ; 
  assign GenStackBus[39].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[39].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[40].mgr__sys__allSynchronized   =  GenStackBus[40].sys__pe__allSynchronized                                ; 
  assign GenStackBus[40].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[40].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[40].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[40].sys__mgr__ready             ; 
  assign GenStackBus[40].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[40].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[41].mgr__sys__allSynchronized   =  GenStackBus[41].sys__pe__allSynchronized                                ; 
  assign GenStackBus[41].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[41].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[41].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[41].sys__mgr__ready             ; 
  assign GenStackBus[41].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[41].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[42].mgr__sys__allSynchronized   =  GenStackBus[42].sys__pe__allSynchronized                                ; 
  assign GenStackBus[42].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[42].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[42].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[42].sys__mgr__ready             ; 
  assign GenStackBus[42].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[42].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[43].mgr__sys__allSynchronized   =  GenStackBus[43].sys__pe__allSynchronized                                ; 
  assign GenStackBus[43].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[43].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[43].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[43].sys__mgr__ready             ; 
  assign GenStackBus[43].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[43].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[44].mgr__sys__allSynchronized   =  GenStackBus[44].sys__pe__allSynchronized                                ; 
  assign GenStackBus[44].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[44].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[44].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[44].sys__mgr__ready             ; 
  assign GenStackBus[44].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[44].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[45].mgr__sys__allSynchronized   =  GenStackBus[45].sys__pe__allSynchronized                                ; 
  assign GenStackBus[45].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[45].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[45].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[45].sys__mgr__ready             ; 
  assign GenStackBus[45].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[45].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[46].mgr__sys__allSynchronized   =  GenStackBus[46].sys__pe__allSynchronized                                ; 
  assign GenStackBus[46].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[46].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[46].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[46].sys__mgr__ready             ; 
  assign GenStackBus[46].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[46].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[47].mgr__sys__allSynchronized   =  GenStackBus[47].sys__pe__allSynchronized                                ; 
  assign GenStackBus[47].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[47].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[47].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[47].sys__mgr__ready             ; 
  assign GenStackBus[47].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[47].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[48].mgr__sys__allSynchronized   =  GenStackBus[48].sys__pe__allSynchronized                                ; 
  assign GenStackBus[48].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[48].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[48].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[48].sys__mgr__ready             ; 
  assign GenStackBus[48].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[48].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[49].mgr__sys__allSynchronized   =  GenStackBus[49].sys__pe__allSynchronized                                ; 
  assign GenStackBus[49].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[49].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[49].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[49].sys__mgr__ready             ; 
  assign GenStackBus[49].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[49].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[50].mgr__sys__allSynchronized   =  GenStackBus[50].sys__pe__allSynchronized                                ; 
  assign GenStackBus[50].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[50].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[50].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[50].sys__mgr__ready             ; 
  assign GenStackBus[50].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[50].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[51].mgr__sys__allSynchronized   =  GenStackBus[51].sys__pe__allSynchronized                                ; 
  assign GenStackBus[51].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[51].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[51].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[51].sys__mgr__ready             ; 
  assign GenStackBus[51].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[51].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[52].mgr__sys__allSynchronized   =  GenStackBus[52].sys__pe__allSynchronized                                ; 
  assign GenStackBus[52].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[52].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[52].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[52].sys__mgr__ready             ; 
  assign GenStackBus[52].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[52].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[53].mgr__sys__allSynchronized   =  GenStackBus[53].sys__pe__allSynchronized                                ; 
  assign GenStackBus[53].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[53].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[53].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[53].sys__mgr__ready             ; 
  assign GenStackBus[53].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[53].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[54].mgr__sys__allSynchronized   =  GenStackBus[54].sys__pe__allSynchronized                                ; 
  assign GenStackBus[54].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[54].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[54].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[54].sys__mgr__ready             ; 
  assign GenStackBus[54].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[54].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[55].mgr__sys__allSynchronized   =  GenStackBus[55].sys__pe__allSynchronized                                ; 
  assign GenStackBus[55].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[55].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[55].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[55].sys__mgr__ready             ; 
  assign GenStackBus[55].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[55].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[56].mgr__sys__allSynchronized   =  GenStackBus[56].sys__pe__allSynchronized                                ; 
  assign GenStackBus[56].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[56].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[56].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[56].sys__mgr__ready             ; 
  assign GenStackBus[56].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[56].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[57].mgr__sys__allSynchronized   =  GenStackBus[57].sys__pe__allSynchronized                                ; 
  assign GenStackBus[57].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[57].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[57].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[57].sys__mgr__ready             ; 
  assign GenStackBus[57].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[57].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[58].mgr__sys__allSynchronized   =  GenStackBus[58].sys__pe__allSynchronized                                ; 
  assign GenStackBus[58].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[58].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[58].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[58].sys__mgr__ready             ; 
  assign GenStackBus[58].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[58].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[59].mgr__sys__allSynchronized   =  GenStackBus[59].sys__pe__allSynchronized                                ; 
  assign GenStackBus[59].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[59].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[59].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[59].sys__mgr__ready             ; 
  assign GenStackBus[59].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[59].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[60].mgr__sys__allSynchronized   =  GenStackBus[60].sys__pe__allSynchronized                                ; 
  assign GenStackBus[60].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[60].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[60].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[60].sys__mgr__ready             ; 
  assign GenStackBus[60].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[60].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[61].mgr__sys__allSynchronized   =  GenStackBus[61].sys__pe__allSynchronized                                ; 
  assign GenStackBus[61].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[61].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[61].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[61].sys__mgr__ready             ; 
  assign GenStackBus[61].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[61].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[62].mgr__sys__allSynchronized   =  GenStackBus[62].sys__pe__allSynchronized                                ; 
  assign GenStackBus[62].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[62].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[62].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[62].sys__mgr__ready             ; 
  assign GenStackBus[62].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[62].sys__mgr__complete          ; 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.   
  assign system_inst.manager_array_inst.mgr_inst[63].mgr__sys__allSynchronized   =  GenStackBus[63].sys__pe__allSynchronized                                ; 
  assign GenStackBus[63].pe__sys__thisSynchronized                               =  system_inst.manager_array_inst.mgr_inst[63].sys__mgr__thisSynchronized  ; 
  assign GenStackBus[63].pe__sys__ready                                          =  system_inst.manager_array_inst.mgr_inst[63].sys__mgr__ready             ; 
  assign GenStackBus[63].pe__sys__complete                                       =  system_inst.manager_array_inst.mgr_inst[63].sys__mgr__complete          ; 
