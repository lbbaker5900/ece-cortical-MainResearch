
//------------------------------------------------
// MEM_ACC_CONT_ARBITER_STATE width
//------------------------------------------------
`define MEM_ACC_CONT_STATE_MSB            68
`define MEM_ACC_CONT_STATE_LSB            0
`define MEM_ACC_CONT_STATE_SIZE           (`MEM_ACC_CONT_STATE_MSB - `MEM_ACC_CONT_STATE_LSB +1)
`define MEM_ACC_CONT_STATE_RANGE           `MEM_ACC_CONT_STATE_MSB : `MEM_ACC_CONT_STATE_LSB

//------------------------------------------------------------------------------------------------
//------------------------------------------------
// MEM_ACC_CONT state machine states
//------------------------------------------------

`define MEM_ACC_CONT_WAIT                    69'd1
`define MEM_ACC_CONT_DMA                     69'd2
`define MEM_ACC_CONT_LDST                    69'd4
`define MEM_ACC_CONT_LDST_READ_ACCESS        69'd8
`define MEM_ACC_CONT_LDST_WRITE_ACCESS       69'd16
`define MEM_ACC_CONT_DMA_STRM0_READ_ACCESS   69'd32
`define MEM_ACC_CONT_DMA_STRM0_WRITE_ACCESS  69'd64
`define MEM_ACC_CONT_DMA_STRM1_READ_ACCESS   69'd128
`define MEM_ACC_CONT_DMA_STRM1_WRITE_ACCESS  69'd256
`define MEM_ACC_CONT_DMA_STRM2_READ_ACCESS   69'd512
`define MEM_ACC_CONT_DMA_STRM2_WRITE_ACCESS  69'd1024
`define MEM_ACC_CONT_DMA_STRM3_READ_ACCESS   69'd2048
`define MEM_ACC_CONT_DMA_STRM3_WRITE_ACCESS  69'd4096
`define MEM_ACC_CONT_DMA_STRM4_READ_ACCESS   69'd8192
`define MEM_ACC_CONT_DMA_STRM4_WRITE_ACCESS  69'd16384
`define MEM_ACC_CONT_DMA_STRM5_READ_ACCESS   69'd32768
`define MEM_ACC_CONT_DMA_STRM5_WRITE_ACCESS  69'd65536
`define MEM_ACC_CONT_DMA_STRM6_READ_ACCESS   69'd131072
`define MEM_ACC_CONT_DMA_STRM6_WRITE_ACCESS  69'd262144
`define MEM_ACC_CONT_DMA_STRM7_READ_ACCESS   69'd524288
`define MEM_ACC_CONT_DMA_STRM7_WRITE_ACCESS  69'd1048576
`define MEM_ACC_CONT_DMA_STRM8_READ_ACCESS   69'd2097152
`define MEM_ACC_CONT_DMA_STRM8_WRITE_ACCESS  69'd4194304
`define MEM_ACC_CONT_DMA_STRM9_READ_ACCESS   69'd8388608
`define MEM_ACC_CONT_DMA_STRM9_WRITE_ACCESS  69'd16777216
`define MEM_ACC_CONT_DMA_STRM10_READ_ACCESS   69'd33554432
`define MEM_ACC_CONT_DMA_STRM10_WRITE_ACCESS  69'd67108864
`define MEM_ACC_CONT_DMA_STRM11_READ_ACCESS   69'd134217728
`define MEM_ACC_CONT_DMA_STRM11_WRITE_ACCESS  69'd268435456
`define MEM_ACC_CONT_DMA_STRM12_READ_ACCESS   69'd536870912
`define MEM_ACC_CONT_DMA_STRM12_WRITE_ACCESS  69'd1073741824
`define MEM_ACC_CONT_DMA_STRM13_READ_ACCESS   69'd2147483648
`define MEM_ACC_CONT_DMA_STRM13_WRITE_ACCESS  69'd4294967296
`define MEM_ACC_CONT_DMA_STRM14_READ_ACCESS   69'd8589934592
`define MEM_ACC_CONT_DMA_STRM14_WRITE_ACCESS  69'd17179869184
`define MEM_ACC_CONT_DMA_STRM15_READ_ACCESS   69'd34359738368
`define MEM_ACC_CONT_DMA_STRM15_WRITE_ACCESS  69'd68719476736
`define MEM_ACC_CONT_DMA_STRM16_READ_ACCESS   69'd137438953472
`define MEM_ACC_CONT_DMA_STRM16_WRITE_ACCESS  69'd274877906944
`define MEM_ACC_CONT_DMA_STRM17_READ_ACCESS   69'd549755813888
`define MEM_ACC_CONT_DMA_STRM17_WRITE_ACCESS  69'd1099511627776
`define MEM_ACC_CONT_DMA_STRM18_READ_ACCESS   69'd2199023255552
`define MEM_ACC_CONT_DMA_STRM18_WRITE_ACCESS  69'd4398046511104
`define MEM_ACC_CONT_DMA_STRM19_READ_ACCESS   69'd8796093022208
`define MEM_ACC_CONT_DMA_STRM19_WRITE_ACCESS  69'd17592186044416
`define MEM_ACC_CONT_DMA_STRM20_READ_ACCESS   69'd35184372088832
`define MEM_ACC_CONT_DMA_STRM20_WRITE_ACCESS  69'd70368744177664
`define MEM_ACC_CONT_DMA_STRM21_READ_ACCESS   69'd140737488355328
`define MEM_ACC_CONT_DMA_STRM21_WRITE_ACCESS  69'd281474976710656
`define MEM_ACC_CONT_DMA_STRM22_READ_ACCESS   69'd562949953421312
`define MEM_ACC_CONT_DMA_STRM22_WRITE_ACCESS  69'd1125899906842624
`define MEM_ACC_CONT_DMA_STRM23_READ_ACCESS   69'd2251799813685248
`define MEM_ACC_CONT_DMA_STRM23_WRITE_ACCESS  69'd4503599627370496
`define MEM_ACC_CONT_DMA_STRM24_READ_ACCESS   69'd9007199254740992
`define MEM_ACC_CONT_DMA_STRM24_WRITE_ACCESS  69'd18014398509481984
`define MEM_ACC_CONT_DMA_STRM25_READ_ACCESS   69'd36028797018963968
`define MEM_ACC_CONT_DMA_STRM25_WRITE_ACCESS  69'd72057594037927936
`define MEM_ACC_CONT_DMA_STRM26_READ_ACCESS   69'd144115188075855872
`define MEM_ACC_CONT_DMA_STRM26_WRITE_ACCESS  69'd288230376151711744
`define MEM_ACC_CONT_DMA_STRM27_READ_ACCESS   69'd576460752303423488
`define MEM_ACC_CONT_DMA_STRM27_WRITE_ACCESS  69'd1152921504606846976
`define MEM_ACC_CONT_DMA_STRM28_READ_ACCESS   69'd2305843009213693952
`define MEM_ACC_CONT_DMA_STRM28_WRITE_ACCESS  69'd4611686018427387904
`define MEM_ACC_CONT_DMA_STRM29_READ_ACCESS   69'd9223372036854775808
`define MEM_ACC_CONT_DMA_STRM29_WRITE_ACCESS  69'd18446744073709551616
`define MEM_ACC_CONT_DMA_STRM30_READ_ACCESS   69'd36893488147419103232
`define MEM_ACC_CONT_DMA_STRM30_WRITE_ACCESS  69'd73786976294838206464
`define MEM_ACC_CONT_DMA_STRM31_READ_ACCESS   69'd147573952589676412928
`define MEM_ACC_CONT_DMA_STRM31_WRITE_ACCESS  69'd295147905179352825856