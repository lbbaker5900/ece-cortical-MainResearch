
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[0].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[0].stu__mgr__valid    ;      
        assign UpstreamStackBus[0].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[0].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[0].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[0].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[0].mgr__stu__ready    ;      
        assign UpstreamStackBus[0].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[0].stu__mgr__type     ;      
        assign UpstreamStackBus[0].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[0].stu__mgr__data     ;      
        assign UpstreamStackBus[0].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[0].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[1].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[1].stu__mgr__valid    ;      
        assign UpstreamStackBus[1].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[1].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[1].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[1].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[1].mgr__stu__ready    ;      
        assign UpstreamStackBus[1].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[1].stu__mgr__type     ;      
        assign UpstreamStackBus[1].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[1].stu__mgr__data     ;      
        assign UpstreamStackBus[1].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[1].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[2].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[2].stu__mgr__valid    ;      
        assign UpstreamStackBus[2].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[2].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[2].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[2].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[2].mgr__stu__ready    ;      
        assign UpstreamStackBus[2].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[2].stu__mgr__type     ;      
        assign UpstreamStackBus[2].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[2].stu__mgr__data     ;      
        assign UpstreamStackBus[2].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[2].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[3].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[3].stu__mgr__valid    ;      
        assign UpstreamStackBus[3].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[3].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[3].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[3].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[3].mgr__stu__ready    ;      
        assign UpstreamStackBus[3].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[3].stu__mgr__type     ;      
        assign UpstreamStackBus[3].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[3].stu__mgr__data     ;      
        assign UpstreamStackBus[3].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[3].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[4].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[4].stu__mgr__valid    ;      
        assign UpstreamStackBus[4].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[4].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[4].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[4].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[4].mgr__stu__ready    ;      
        assign UpstreamStackBus[4].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[4].stu__mgr__type     ;      
        assign UpstreamStackBus[4].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[4].stu__mgr__data     ;      
        assign UpstreamStackBus[4].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[4].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[5].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[5].stu__mgr__valid    ;      
        assign UpstreamStackBus[5].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[5].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[5].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[5].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[5].mgr__stu__ready    ;      
        assign UpstreamStackBus[5].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[5].stu__mgr__type     ;      
        assign UpstreamStackBus[5].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[5].stu__mgr__data     ;      
        assign UpstreamStackBus[5].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[5].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[6].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[6].stu__mgr__valid    ;      
        assign UpstreamStackBus[6].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[6].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[6].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[6].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[6].mgr__stu__ready    ;      
        assign UpstreamStackBus[6].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[6].stu__mgr__type     ;      
        assign UpstreamStackBus[6].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[6].stu__mgr__data     ;      
        assign UpstreamStackBus[6].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[6].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[7].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[7].stu__mgr__valid    ;      
        assign UpstreamStackBus[7].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[7].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[7].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[7].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[7].mgr__stu__ready    ;      
        assign UpstreamStackBus[7].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[7].stu__mgr__type     ;      
        assign UpstreamStackBus[7].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[7].stu__mgr__data     ;      
        assign UpstreamStackBus[7].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[7].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[8].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[8].stu__mgr__valid    ;      
        assign UpstreamStackBus[8].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[8].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[8].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[8].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[8].mgr__stu__ready    ;      
        assign UpstreamStackBus[8].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[8].stu__mgr__type     ;      
        assign UpstreamStackBus[8].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[8].stu__mgr__data     ;      
        assign UpstreamStackBus[8].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[8].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[9].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[9].stu__mgr__valid    ;      
        assign UpstreamStackBus[9].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[9].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[9].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[9].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[9].mgr__stu__ready    ;      
        assign UpstreamStackBus[9].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[9].stu__mgr__type     ;      
        assign UpstreamStackBus[9].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[9].stu__mgr__data     ;      
        assign UpstreamStackBus[9].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[9].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[10].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[10].stu__mgr__valid    ;      
        assign UpstreamStackBus[10].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[10].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[10].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[10].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[10].mgr__stu__ready    ;      
        assign UpstreamStackBus[10].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[10].stu__mgr__type     ;      
        assign UpstreamStackBus[10].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[10].stu__mgr__data     ;      
        assign UpstreamStackBus[10].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[10].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[11].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[11].stu__mgr__valid    ;      
        assign UpstreamStackBus[11].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[11].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[11].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[11].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[11].mgr__stu__ready    ;      
        assign UpstreamStackBus[11].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[11].stu__mgr__type     ;      
        assign UpstreamStackBus[11].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[11].stu__mgr__data     ;      
        assign UpstreamStackBus[11].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[11].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[12].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[12].stu__mgr__valid    ;      
        assign UpstreamStackBus[12].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[12].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[12].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[12].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[12].mgr__stu__ready    ;      
        assign UpstreamStackBus[12].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[12].stu__mgr__type     ;      
        assign UpstreamStackBus[12].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[12].stu__mgr__data     ;      
        assign UpstreamStackBus[12].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[12].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[13].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[13].stu__mgr__valid    ;      
        assign UpstreamStackBus[13].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[13].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[13].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[13].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[13].mgr__stu__ready    ;      
        assign UpstreamStackBus[13].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[13].stu__mgr__type     ;      
        assign UpstreamStackBus[13].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[13].stu__mgr__data     ;      
        assign UpstreamStackBus[13].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[13].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[14].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[14].stu__mgr__valid    ;      
        assign UpstreamStackBus[14].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[14].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[14].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[14].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[14].mgr__stu__ready    ;      
        assign UpstreamStackBus[14].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[14].stu__mgr__type     ;      
        assign UpstreamStackBus[14].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[14].stu__mgr__data     ;      
        assign UpstreamStackBus[14].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[14].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[15].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[15].stu__mgr__valid    ;      
        assign UpstreamStackBus[15].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[15].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[15].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[15].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[15].mgr__stu__ready    ;      
        assign UpstreamStackBus[15].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[15].stu__mgr__type     ;      
        assign UpstreamStackBus[15].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[15].stu__mgr__data     ;      
        assign UpstreamStackBus[15].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[15].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[16].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[16].stu__mgr__valid    ;      
        assign UpstreamStackBus[16].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[16].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[16].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[16].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[16].mgr__stu__ready    ;      
        assign UpstreamStackBus[16].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[16].stu__mgr__type     ;      
        assign UpstreamStackBus[16].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[16].stu__mgr__data     ;      
        assign UpstreamStackBus[16].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[16].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[17].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[17].stu__mgr__valid    ;      
        assign UpstreamStackBus[17].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[17].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[17].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[17].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[17].mgr__stu__ready    ;      
        assign UpstreamStackBus[17].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[17].stu__mgr__type     ;      
        assign UpstreamStackBus[17].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[17].stu__mgr__data     ;      
        assign UpstreamStackBus[17].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[17].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[18].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[18].stu__mgr__valid    ;      
        assign UpstreamStackBus[18].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[18].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[18].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[18].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[18].mgr__stu__ready    ;      
        assign UpstreamStackBus[18].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[18].stu__mgr__type     ;      
        assign UpstreamStackBus[18].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[18].stu__mgr__data     ;      
        assign UpstreamStackBus[18].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[18].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[19].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[19].stu__mgr__valid    ;      
        assign UpstreamStackBus[19].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[19].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[19].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[19].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[19].mgr__stu__ready    ;      
        assign UpstreamStackBus[19].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[19].stu__mgr__type     ;      
        assign UpstreamStackBus[19].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[19].stu__mgr__data     ;      
        assign UpstreamStackBus[19].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[19].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[20].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[20].stu__mgr__valid    ;      
        assign UpstreamStackBus[20].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[20].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[20].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[20].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[20].mgr__stu__ready    ;      
        assign UpstreamStackBus[20].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[20].stu__mgr__type     ;      
        assign UpstreamStackBus[20].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[20].stu__mgr__data     ;      
        assign UpstreamStackBus[20].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[20].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[21].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[21].stu__mgr__valid    ;      
        assign UpstreamStackBus[21].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[21].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[21].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[21].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[21].mgr__stu__ready    ;      
        assign UpstreamStackBus[21].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[21].stu__mgr__type     ;      
        assign UpstreamStackBus[21].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[21].stu__mgr__data     ;      
        assign UpstreamStackBus[21].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[21].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[22].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[22].stu__mgr__valid    ;      
        assign UpstreamStackBus[22].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[22].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[22].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[22].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[22].mgr__stu__ready    ;      
        assign UpstreamStackBus[22].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[22].stu__mgr__type     ;      
        assign UpstreamStackBus[22].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[22].stu__mgr__data     ;      
        assign UpstreamStackBus[22].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[22].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[23].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[23].stu__mgr__valid    ;      
        assign UpstreamStackBus[23].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[23].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[23].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[23].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[23].mgr__stu__ready    ;      
        assign UpstreamStackBus[23].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[23].stu__mgr__type     ;      
        assign UpstreamStackBus[23].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[23].stu__mgr__data     ;      
        assign UpstreamStackBus[23].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[23].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[24].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[24].stu__mgr__valid    ;      
        assign UpstreamStackBus[24].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[24].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[24].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[24].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[24].mgr__stu__ready    ;      
        assign UpstreamStackBus[24].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[24].stu__mgr__type     ;      
        assign UpstreamStackBus[24].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[24].stu__mgr__data     ;      
        assign UpstreamStackBus[24].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[24].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[25].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[25].stu__mgr__valid    ;      
        assign UpstreamStackBus[25].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[25].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[25].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[25].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[25].mgr__stu__ready    ;      
        assign UpstreamStackBus[25].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[25].stu__mgr__type     ;      
        assign UpstreamStackBus[25].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[25].stu__mgr__data     ;      
        assign UpstreamStackBus[25].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[25].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[26].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[26].stu__mgr__valid    ;      
        assign UpstreamStackBus[26].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[26].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[26].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[26].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[26].mgr__stu__ready    ;      
        assign UpstreamStackBus[26].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[26].stu__mgr__type     ;      
        assign UpstreamStackBus[26].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[26].stu__mgr__data     ;      
        assign UpstreamStackBus[26].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[26].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[27].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[27].stu__mgr__valid    ;      
        assign UpstreamStackBus[27].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[27].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[27].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[27].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[27].mgr__stu__ready    ;      
        assign UpstreamStackBus[27].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[27].stu__mgr__type     ;      
        assign UpstreamStackBus[27].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[27].stu__mgr__data     ;      
        assign UpstreamStackBus[27].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[27].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[28].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[28].stu__mgr__valid    ;      
        assign UpstreamStackBus[28].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[28].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[28].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[28].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[28].mgr__stu__ready    ;      
        assign UpstreamStackBus[28].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[28].stu__mgr__type     ;      
        assign UpstreamStackBus[28].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[28].stu__mgr__data     ;      
        assign UpstreamStackBus[28].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[28].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[29].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[29].stu__mgr__valid    ;      
        assign UpstreamStackBus[29].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[29].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[29].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[29].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[29].mgr__stu__ready    ;      
        assign UpstreamStackBus[29].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[29].stu__mgr__type     ;      
        assign UpstreamStackBus[29].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[29].stu__mgr__data     ;      
        assign UpstreamStackBus[29].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[29].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[30].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[30].stu__mgr__valid    ;      
        assign UpstreamStackBus[30].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[30].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[30].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[30].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[30].mgr__stu__ready    ;      
        assign UpstreamStackBus[30].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[30].stu__mgr__type     ;      
        assign UpstreamStackBus[30].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[30].stu__mgr__data     ;      
        assign UpstreamStackBus[30].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[30].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[31].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[31].stu__mgr__valid    ;      
        assign UpstreamStackBus[31].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[31].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[31].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[31].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[31].mgr__stu__ready    ;      
        assign UpstreamStackBus[31].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[31].stu__mgr__type     ;      
        assign UpstreamStackBus[31].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[31].stu__mgr__data     ;      
        assign UpstreamStackBus[31].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[31].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[32].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[32].stu__mgr__valid    ;      
        assign UpstreamStackBus[32].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[32].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[32].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[32].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[32].mgr__stu__ready    ;      
        assign UpstreamStackBus[32].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[32].stu__mgr__type     ;      
        assign UpstreamStackBus[32].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[32].stu__mgr__data     ;      
        assign UpstreamStackBus[32].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[32].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[33].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[33].stu__mgr__valid    ;      
        assign UpstreamStackBus[33].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[33].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[33].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[33].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[33].mgr__stu__ready    ;      
        assign UpstreamStackBus[33].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[33].stu__mgr__type     ;      
        assign UpstreamStackBus[33].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[33].stu__mgr__data     ;      
        assign UpstreamStackBus[33].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[33].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[34].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[34].stu__mgr__valid    ;      
        assign UpstreamStackBus[34].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[34].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[34].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[34].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[34].mgr__stu__ready    ;      
        assign UpstreamStackBus[34].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[34].stu__mgr__type     ;      
        assign UpstreamStackBus[34].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[34].stu__mgr__data     ;      
        assign UpstreamStackBus[34].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[34].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[35].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[35].stu__mgr__valid    ;      
        assign UpstreamStackBus[35].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[35].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[35].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[35].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[35].mgr__stu__ready    ;      
        assign UpstreamStackBus[35].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[35].stu__mgr__type     ;      
        assign UpstreamStackBus[35].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[35].stu__mgr__data     ;      
        assign UpstreamStackBus[35].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[35].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[36].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[36].stu__mgr__valid    ;      
        assign UpstreamStackBus[36].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[36].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[36].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[36].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[36].mgr__stu__ready    ;      
        assign UpstreamStackBus[36].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[36].stu__mgr__type     ;      
        assign UpstreamStackBus[36].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[36].stu__mgr__data     ;      
        assign UpstreamStackBus[36].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[36].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[37].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[37].stu__mgr__valid    ;      
        assign UpstreamStackBus[37].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[37].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[37].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[37].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[37].mgr__stu__ready    ;      
        assign UpstreamStackBus[37].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[37].stu__mgr__type     ;      
        assign UpstreamStackBus[37].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[37].stu__mgr__data     ;      
        assign UpstreamStackBus[37].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[37].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[38].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[38].stu__mgr__valid    ;      
        assign UpstreamStackBus[38].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[38].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[38].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[38].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[38].mgr__stu__ready    ;      
        assign UpstreamStackBus[38].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[38].stu__mgr__type     ;      
        assign UpstreamStackBus[38].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[38].stu__mgr__data     ;      
        assign UpstreamStackBus[38].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[38].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[39].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[39].stu__mgr__valid    ;      
        assign UpstreamStackBus[39].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[39].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[39].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[39].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[39].mgr__stu__ready    ;      
        assign UpstreamStackBus[39].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[39].stu__mgr__type     ;      
        assign UpstreamStackBus[39].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[39].stu__mgr__data     ;      
        assign UpstreamStackBus[39].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[39].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[40].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[40].stu__mgr__valid    ;      
        assign UpstreamStackBus[40].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[40].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[40].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[40].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[40].mgr__stu__ready    ;      
        assign UpstreamStackBus[40].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[40].stu__mgr__type     ;      
        assign UpstreamStackBus[40].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[40].stu__mgr__data     ;      
        assign UpstreamStackBus[40].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[40].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[41].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[41].stu__mgr__valid    ;      
        assign UpstreamStackBus[41].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[41].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[41].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[41].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[41].mgr__stu__ready    ;      
        assign UpstreamStackBus[41].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[41].stu__mgr__type     ;      
        assign UpstreamStackBus[41].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[41].stu__mgr__data     ;      
        assign UpstreamStackBus[41].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[41].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[42].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[42].stu__mgr__valid    ;      
        assign UpstreamStackBus[42].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[42].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[42].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[42].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[42].mgr__stu__ready    ;      
        assign UpstreamStackBus[42].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[42].stu__mgr__type     ;      
        assign UpstreamStackBus[42].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[42].stu__mgr__data     ;      
        assign UpstreamStackBus[42].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[42].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[43].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[43].stu__mgr__valid    ;      
        assign UpstreamStackBus[43].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[43].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[43].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[43].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[43].mgr__stu__ready    ;      
        assign UpstreamStackBus[43].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[43].stu__mgr__type     ;      
        assign UpstreamStackBus[43].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[43].stu__mgr__data     ;      
        assign UpstreamStackBus[43].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[43].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[44].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[44].stu__mgr__valid    ;      
        assign UpstreamStackBus[44].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[44].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[44].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[44].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[44].mgr__stu__ready    ;      
        assign UpstreamStackBus[44].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[44].stu__mgr__type     ;      
        assign UpstreamStackBus[44].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[44].stu__mgr__data     ;      
        assign UpstreamStackBus[44].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[44].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[45].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[45].stu__mgr__valid    ;      
        assign UpstreamStackBus[45].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[45].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[45].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[45].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[45].mgr__stu__ready    ;      
        assign UpstreamStackBus[45].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[45].stu__mgr__type     ;      
        assign UpstreamStackBus[45].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[45].stu__mgr__data     ;      
        assign UpstreamStackBus[45].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[45].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[46].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[46].stu__mgr__valid    ;      
        assign UpstreamStackBus[46].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[46].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[46].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[46].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[46].mgr__stu__ready    ;      
        assign UpstreamStackBus[46].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[46].stu__mgr__type     ;      
        assign UpstreamStackBus[46].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[46].stu__mgr__data     ;      
        assign UpstreamStackBus[46].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[46].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[47].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[47].stu__mgr__valid    ;      
        assign UpstreamStackBus[47].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[47].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[47].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[47].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[47].mgr__stu__ready    ;      
        assign UpstreamStackBus[47].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[47].stu__mgr__type     ;      
        assign UpstreamStackBus[47].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[47].stu__mgr__data     ;      
        assign UpstreamStackBus[47].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[47].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[48].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[48].stu__mgr__valid    ;      
        assign UpstreamStackBus[48].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[48].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[48].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[48].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[48].mgr__stu__ready    ;      
        assign UpstreamStackBus[48].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[48].stu__mgr__type     ;      
        assign UpstreamStackBus[48].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[48].stu__mgr__data     ;      
        assign UpstreamStackBus[48].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[48].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[49].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[49].stu__mgr__valid    ;      
        assign UpstreamStackBus[49].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[49].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[49].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[49].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[49].mgr__stu__ready    ;      
        assign UpstreamStackBus[49].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[49].stu__mgr__type     ;      
        assign UpstreamStackBus[49].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[49].stu__mgr__data     ;      
        assign UpstreamStackBus[49].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[49].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[50].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[50].stu__mgr__valid    ;      
        assign UpstreamStackBus[50].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[50].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[50].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[50].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[50].mgr__stu__ready    ;      
        assign UpstreamStackBus[50].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[50].stu__mgr__type     ;      
        assign UpstreamStackBus[50].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[50].stu__mgr__data     ;      
        assign UpstreamStackBus[50].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[50].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[51].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[51].stu__mgr__valid    ;      
        assign UpstreamStackBus[51].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[51].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[51].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[51].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[51].mgr__stu__ready    ;      
        assign UpstreamStackBus[51].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[51].stu__mgr__type     ;      
        assign UpstreamStackBus[51].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[51].stu__mgr__data     ;      
        assign UpstreamStackBus[51].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[51].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[52].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[52].stu__mgr__valid    ;      
        assign UpstreamStackBus[52].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[52].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[52].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[52].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[52].mgr__stu__ready    ;      
        assign UpstreamStackBus[52].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[52].stu__mgr__type     ;      
        assign UpstreamStackBus[52].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[52].stu__mgr__data     ;      
        assign UpstreamStackBus[52].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[52].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[53].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[53].stu__mgr__valid    ;      
        assign UpstreamStackBus[53].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[53].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[53].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[53].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[53].mgr__stu__ready    ;      
        assign UpstreamStackBus[53].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[53].stu__mgr__type     ;      
        assign UpstreamStackBus[53].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[53].stu__mgr__data     ;      
        assign UpstreamStackBus[53].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[53].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[54].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[54].stu__mgr__valid    ;      
        assign UpstreamStackBus[54].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[54].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[54].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[54].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[54].mgr__stu__ready    ;      
        assign UpstreamStackBus[54].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[54].stu__mgr__type     ;      
        assign UpstreamStackBus[54].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[54].stu__mgr__data     ;      
        assign UpstreamStackBus[54].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[54].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[55].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[55].stu__mgr__valid    ;      
        assign UpstreamStackBus[55].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[55].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[55].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[55].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[55].mgr__stu__ready    ;      
        assign UpstreamStackBus[55].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[55].stu__mgr__type     ;      
        assign UpstreamStackBus[55].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[55].stu__mgr__data     ;      
        assign UpstreamStackBus[55].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[55].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[56].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[56].stu__mgr__valid    ;      
        assign UpstreamStackBus[56].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[56].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[56].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[56].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[56].mgr__stu__ready    ;      
        assign UpstreamStackBus[56].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[56].stu__mgr__type     ;      
        assign UpstreamStackBus[56].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[56].stu__mgr__data     ;      
        assign UpstreamStackBus[56].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[56].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[57].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[57].stu__mgr__valid    ;      
        assign UpstreamStackBus[57].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[57].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[57].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[57].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[57].mgr__stu__ready    ;      
        assign UpstreamStackBus[57].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[57].stu__mgr__type     ;      
        assign UpstreamStackBus[57].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[57].stu__mgr__data     ;      
        assign UpstreamStackBus[57].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[57].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[58].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[58].stu__mgr__valid    ;      
        assign UpstreamStackBus[58].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[58].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[58].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[58].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[58].mgr__stu__ready    ;      
        assign UpstreamStackBus[58].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[58].stu__mgr__type     ;      
        assign UpstreamStackBus[58].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[58].stu__mgr__data     ;      
        assign UpstreamStackBus[58].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[58].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[59].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[59].stu__mgr__valid    ;      
        assign UpstreamStackBus[59].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[59].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[59].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[59].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[59].mgr__stu__ready    ;      
        assign UpstreamStackBus[59].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[59].stu__mgr__type     ;      
        assign UpstreamStackBus[59].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[59].stu__mgr__data     ;      
        assign UpstreamStackBus[59].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[59].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[60].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[60].stu__mgr__valid    ;      
        assign UpstreamStackBus[60].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[60].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[60].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[60].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[60].mgr__stu__ready    ;      
        assign UpstreamStackBus[60].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[60].stu__mgr__type     ;      
        assign UpstreamStackBus[60].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[60].stu__mgr__data     ;      
        assign UpstreamStackBus[60].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[60].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[61].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[61].stu__mgr__valid    ;      
        assign UpstreamStackBus[61].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[61].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[61].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[61].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[61].mgr__stu__ready    ;      
        assign UpstreamStackBus[61].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[61].stu__mgr__type     ;      
        assign UpstreamStackBus[61].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[61].stu__mgr__data     ;      
        assign UpstreamStackBus[61].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[61].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[62].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[62].stu__mgr__valid    ;      
        assign UpstreamStackBus[62].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[62].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[62].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[62].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[62].mgr__stu__ready    ;      
        assign UpstreamStackBus[62].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[62].stu__mgr__type     ;      
        assign UpstreamStackBus[62].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[62].stu__mgr__data     ;      
        assign UpstreamStackBus[62].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[62].stu__mgr__oob_data ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign UpstreamStackBus[63].pe__stu__valid                                =   system_inst.manager_array_inst.mgr_inst[63].stu__mgr__valid    ;      
        assign UpstreamStackBus[63].pe__stu__cntl                                 =   system_inst.manager_array_inst.mgr_inst[63].stu__mgr__cntl     ;      
        // manager module stu_cntl now driving ready, so just capture state of ready                                                                                                          
        //assign system_inst.manager_array_inst.mgr_inst[63].mgr__stu__ready        =   1'b1                                                           ;      
        assign UpstreamStackBus[63].stu__pe__ready                                =   system_inst.manager_array_inst.mgr_inst[63].mgr__stu__ready    ;      
        assign UpstreamStackBus[63].pe__stu__type                                 =   system_inst.manager_array_inst.mgr_inst[63].stu__mgr__type     ;      
        assign UpstreamStackBus[63].pe__stu__data                                 =   system_inst.manager_array_inst.mgr_inst[63].stu__mgr__data     ;      
        assign UpstreamStackBus[63].pe__stu__oob_data                             =   system_inst.manager_array_inst.mgr_inst[63].stu__mgr__oob_data ;      
        