
    // MGR0, Port0 next hop mask                 
    assign mgr_inst[0].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR0_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR0, Port1 next hop mask                 
    assign mgr_inst[0].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR0_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR0, Port2 next hop mask                 
    assign mgr_inst[0].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR0_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR0, Port3 next hop mask                 
    assign mgr_inst[0].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR0_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR1, Port0 next hop mask                 
    assign mgr_inst[1].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR1_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR1, Port1 next hop mask                 
    assign mgr_inst[1].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR1_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR1, Port2 next hop mask                 
    assign mgr_inst[1].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR1_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR1, Port3 next hop mask                 
    assign mgr_inst[1].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR1_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR2, Port0 next hop mask                 
    assign mgr_inst[2].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR2_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR2, Port1 next hop mask                 
    assign mgr_inst[2].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR2_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR2, Port2 next hop mask                 
    assign mgr_inst[2].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR2_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR2, Port3 next hop mask                 
    assign mgr_inst[2].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR2_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR3, Port0 next hop mask                 
    assign mgr_inst[3].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR3_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR3, Port1 next hop mask                 
    assign mgr_inst[3].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR3_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR3, Port2 next hop mask                 
    assign mgr_inst[3].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR3_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR3, Port3 next hop mask                 
    assign mgr_inst[3].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR3_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR4, Port0 next hop mask                 
    assign mgr_inst[4].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR4_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR4, Port1 next hop mask                 
    assign mgr_inst[4].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR4_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR4, Port2 next hop mask                 
    assign mgr_inst[4].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR4_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR4, Port3 next hop mask                 
    assign mgr_inst[4].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR4_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR5, Port0 next hop mask                 
    assign mgr_inst[5].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR5_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR5, Port1 next hop mask                 
    assign mgr_inst[5].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR5_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR5, Port2 next hop mask                 
    assign mgr_inst[5].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR5_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR5, Port3 next hop mask                 
    assign mgr_inst[5].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR5_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR6, Port0 next hop mask                 
    assign mgr_inst[6].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR6_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR6, Port1 next hop mask                 
    assign mgr_inst[6].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR6_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR6, Port2 next hop mask                 
    assign mgr_inst[6].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR6_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR6, Port3 next hop mask                 
    assign mgr_inst[6].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR6_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR7, Port0 next hop mask                 
    assign mgr_inst[7].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR7_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR7, Port1 next hop mask                 
    assign mgr_inst[7].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR7_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR7, Port2 next hop mask                 
    assign mgr_inst[7].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR7_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR7, Port3 next hop mask                 
    assign mgr_inst[7].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR7_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR8, Port0 next hop mask                 
    assign mgr_inst[8].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR8_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR8, Port1 next hop mask                 
    assign mgr_inst[8].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR8_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR8, Port2 next hop mask                 
    assign mgr_inst[8].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR8_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR8, Port3 next hop mask                 
    assign mgr_inst[8].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR8_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR9, Port0 next hop mask                 
    assign mgr_inst[9].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR9_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR9, Port1 next hop mask                 
    assign mgr_inst[9].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR9_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR9, Port2 next hop mask                 
    assign mgr_inst[9].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR9_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR9, Port3 next hop mask                 
    assign mgr_inst[9].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR9_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR10, Port0 next hop mask                 
    assign mgr_inst[10].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR10_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR10, Port1 next hop mask                 
    assign mgr_inst[10].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR10_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR10, Port2 next hop mask                 
    assign mgr_inst[10].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR10_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR10, Port3 next hop mask                 
    assign mgr_inst[10].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR10_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR11, Port0 next hop mask                 
    assign mgr_inst[11].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR11_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR11, Port1 next hop mask                 
    assign mgr_inst[11].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR11_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR11, Port2 next hop mask                 
    assign mgr_inst[11].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR11_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR11, Port3 next hop mask                 
    assign mgr_inst[11].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR11_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR12, Port0 next hop mask                 
    assign mgr_inst[12].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR12_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR12, Port1 next hop mask                 
    assign mgr_inst[12].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR12_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR12, Port2 next hop mask                 
    assign mgr_inst[12].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR12_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR12, Port3 next hop mask                 
    assign mgr_inst[12].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR12_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR13, Port0 next hop mask                 
    assign mgr_inst[13].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR13_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR13, Port1 next hop mask                 
    assign mgr_inst[13].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR13_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR13, Port2 next hop mask                 
    assign mgr_inst[13].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR13_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR13, Port3 next hop mask                 
    assign mgr_inst[13].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR13_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR14, Port0 next hop mask                 
    assign mgr_inst[14].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR14_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR14, Port1 next hop mask                 
    assign mgr_inst[14].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR14_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR14, Port2 next hop mask                 
    assign mgr_inst[14].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR14_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR14, Port3 next hop mask                 
    assign mgr_inst[14].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR14_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR15, Port0 next hop mask                 
    assign mgr_inst[15].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR15_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR15, Port1 next hop mask                 
    assign mgr_inst[15].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR15_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR15, Port2 next hop mask                 
    assign mgr_inst[15].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR15_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR15, Port3 next hop mask                 
    assign mgr_inst[15].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR15_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR16, Port0 next hop mask                 
    assign mgr_inst[16].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR16_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR16, Port1 next hop mask                 
    assign mgr_inst[16].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR16_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR16, Port2 next hop mask                 
    assign mgr_inst[16].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR16_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR16, Port3 next hop mask                 
    assign mgr_inst[16].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR16_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR17, Port0 next hop mask                 
    assign mgr_inst[17].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR17_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR17, Port1 next hop mask                 
    assign mgr_inst[17].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR17_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR17, Port2 next hop mask                 
    assign mgr_inst[17].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR17_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR17, Port3 next hop mask                 
    assign mgr_inst[17].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR17_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR18, Port0 next hop mask                 
    assign mgr_inst[18].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR18_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR18, Port1 next hop mask                 
    assign mgr_inst[18].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR18_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR18, Port2 next hop mask                 
    assign mgr_inst[18].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR18_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR18, Port3 next hop mask                 
    assign mgr_inst[18].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR18_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR19, Port0 next hop mask                 
    assign mgr_inst[19].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR19_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR19, Port1 next hop mask                 
    assign mgr_inst[19].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR19_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR19, Port2 next hop mask                 
    assign mgr_inst[19].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR19_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR19, Port3 next hop mask                 
    assign mgr_inst[19].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR19_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR20, Port0 next hop mask                 
    assign mgr_inst[20].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR20_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR20, Port1 next hop mask                 
    assign mgr_inst[20].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR20_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR20, Port2 next hop mask                 
    assign mgr_inst[20].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR20_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR20, Port3 next hop mask                 
    assign mgr_inst[20].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR20_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR21, Port0 next hop mask                 
    assign mgr_inst[21].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR21_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR21, Port1 next hop mask                 
    assign mgr_inst[21].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR21_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR21, Port2 next hop mask                 
    assign mgr_inst[21].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR21_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR21, Port3 next hop mask                 
    assign mgr_inst[21].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR21_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR22, Port0 next hop mask                 
    assign mgr_inst[22].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR22_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR22, Port1 next hop mask                 
    assign mgr_inst[22].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR22_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR22, Port2 next hop mask                 
    assign mgr_inst[22].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR22_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR22, Port3 next hop mask                 
    assign mgr_inst[22].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR22_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR23, Port0 next hop mask                 
    assign mgr_inst[23].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR23_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR23, Port1 next hop mask                 
    assign mgr_inst[23].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR23_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR23, Port2 next hop mask                 
    assign mgr_inst[23].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR23_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR23, Port3 next hop mask                 
    assign mgr_inst[23].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR23_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR24, Port0 next hop mask                 
    assign mgr_inst[24].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR24_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR24, Port1 next hop mask                 
    assign mgr_inst[24].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR24_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR24, Port2 next hop mask                 
    assign mgr_inst[24].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR24_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR24, Port3 next hop mask                 
    assign mgr_inst[24].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR24_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR25, Port0 next hop mask                 
    assign mgr_inst[25].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR25_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR25, Port1 next hop mask                 
    assign mgr_inst[25].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR25_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR25, Port2 next hop mask                 
    assign mgr_inst[25].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR25_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR25, Port3 next hop mask                 
    assign mgr_inst[25].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR25_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR26, Port0 next hop mask                 
    assign mgr_inst[26].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR26_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR26, Port1 next hop mask                 
    assign mgr_inst[26].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR26_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR26, Port2 next hop mask                 
    assign mgr_inst[26].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR26_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR26, Port3 next hop mask                 
    assign mgr_inst[26].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR26_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR27, Port0 next hop mask                 
    assign mgr_inst[27].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR27_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR27, Port1 next hop mask                 
    assign mgr_inst[27].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR27_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR27, Port2 next hop mask                 
    assign mgr_inst[27].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR27_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR27, Port3 next hop mask                 
    assign mgr_inst[27].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR27_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR28, Port0 next hop mask                 
    assign mgr_inst[28].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR28_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR28, Port1 next hop mask                 
    assign mgr_inst[28].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR28_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR28, Port2 next hop mask                 
    assign mgr_inst[28].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR28_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR28, Port3 next hop mask                 
    assign mgr_inst[28].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR28_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR29, Port0 next hop mask                 
    assign mgr_inst[29].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR29_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR29, Port1 next hop mask                 
    assign mgr_inst[29].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR29_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR29, Port2 next hop mask                 
    assign mgr_inst[29].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR29_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR29, Port3 next hop mask                 
    assign mgr_inst[29].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR29_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR30, Port0 next hop mask                 
    assign mgr_inst[30].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR30_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR30, Port1 next hop mask                 
    assign mgr_inst[30].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR30_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR30, Port2 next hop mask                 
    assign mgr_inst[30].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR30_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR30, Port3 next hop mask                 
    assign mgr_inst[30].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR30_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR31, Port0 next hop mask                 
    assign mgr_inst[31].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR31_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR31, Port1 next hop mask                 
    assign mgr_inst[31].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR31_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR31, Port2 next hop mask                 
    assign mgr_inst[31].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR31_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR31, Port3 next hop mask                 
    assign mgr_inst[31].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR31_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR32, Port0 next hop mask                 
    assign mgr_inst[32].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR32_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR32, Port1 next hop mask                 
    assign mgr_inst[32].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR32_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR32, Port2 next hop mask                 
    assign mgr_inst[32].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR32_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR32, Port3 next hop mask                 
    assign mgr_inst[32].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR32_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR33, Port0 next hop mask                 
    assign mgr_inst[33].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR33_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR33, Port1 next hop mask                 
    assign mgr_inst[33].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR33_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR33, Port2 next hop mask                 
    assign mgr_inst[33].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR33_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR33, Port3 next hop mask                 
    assign mgr_inst[33].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR33_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR34, Port0 next hop mask                 
    assign mgr_inst[34].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR34_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR34, Port1 next hop mask                 
    assign mgr_inst[34].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR34_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR34, Port2 next hop mask                 
    assign mgr_inst[34].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR34_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR34, Port3 next hop mask                 
    assign mgr_inst[34].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR34_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR35, Port0 next hop mask                 
    assign mgr_inst[35].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR35_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR35, Port1 next hop mask                 
    assign mgr_inst[35].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR35_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR35, Port2 next hop mask                 
    assign mgr_inst[35].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR35_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR35, Port3 next hop mask                 
    assign mgr_inst[35].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR35_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR36, Port0 next hop mask                 
    assign mgr_inst[36].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR36_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR36, Port1 next hop mask                 
    assign mgr_inst[36].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR36_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR36, Port2 next hop mask                 
    assign mgr_inst[36].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR36_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR36, Port3 next hop mask                 
    assign mgr_inst[36].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR36_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR37, Port0 next hop mask                 
    assign mgr_inst[37].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR37_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR37, Port1 next hop mask                 
    assign mgr_inst[37].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR37_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR37, Port2 next hop mask                 
    assign mgr_inst[37].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR37_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR37, Port3 next hop mask                 
    assign mgr_inst[37].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR37_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR38, Port0 next hop mask                 
    assign mgr_inst[38].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR38_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR38, Port1 next hop mask                 
    assign mgr_inst[38].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR38_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR38, Port2 next hop mask                 
    assign mgr_inst[38].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR38_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR38, Port3 next hop mask                 
    assign mgr_inst[38].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR38_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR39, Port0 next hop mask                 
    assign mgr_inst[39].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR39_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR39, Port1 next hop mask                 
    assign mgr_inst[39].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR39_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR39, Port2 next hop mask                 
    assign mgr_inst[39].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR39_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR39, Port3 next hop mask                 
    assign mgr_inst[39].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR39_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR40, Port0 next hop mask                 
    assign mgr_inst[40].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR40_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR40, Port1 next hop mask                 
    assign mgr_inst[40].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR40_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR40, Port2 next hop mask                 
    assign mgr_inst[40].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR40_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR40, Port3 next hop mask                 
    assign mgr_inst[40].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR40_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR41, Port0 next hop mask                 
    assign mgr_inst[41].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR41_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR41, Port1 next hop mask                 
    assign mgr_inst[41].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR41_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR41, Port2 next hop mask                 
    assign mgr_inst[41].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR41_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR41, Port3 next hop mask                 
    assign mgr_inst[41].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR41_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR42, Port0 next hop mask                 
    assign mgr_inst[42].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR42_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR42, Port1 next hop mask                 
    assign mgr_inst[42].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR42_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR42, Port2 next hop mask                 
    assign mgr_inst[42].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR42_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR42, Port3 next hop mask                 
    assign mgr_inst[42].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR42_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR43, Port0 next hop mask                 
    assign mgr_inst[43].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR43_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR43, Port1 next hop mask                 
    assign mgr_inst[43].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR43_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR43, Port2 next hop mask                 
    assign mgr_inst[43].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR43_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR43, Port3 next hop mask                 
    assign mgr_inst[43].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR43_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR44, Port0 next hop mask                 
    assign mgr_inst[44].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR44_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR44, Port1 next hop mask                 
    assign mgr_inst[44].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR44_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR44, Port2 next hop mask                 
    assign mgr_inst[44].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR44_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR44, Port3 next hop mask                 
    assign mgr_inst[44].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR44_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR45, Port0 next hop mask                 
    assign mgr_inst[45].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR45_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR45, Port1 next hop mask                 
    assign mgr_inst[45].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR45_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR45, Port2 next hop mask                 
    assign mgr_inst[45].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR45_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR45, Port3 next hop mask                 
    assign mgr_inst[45].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR45_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR46, Port0 next hop mask                 
    assign mgr_inst[46].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR46_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR46, Port1 next hop mask                 
    assign mgr_inst[46].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR46_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR46, Port2 next hop mask                 
    assign mgr_inst[46].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR46_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR46, Port3 next hop mask                 
    assign mgr_inst[46].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR46_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR47, Port0 next hop mask                 
    assign mgr_inst[47].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR47_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR47, Port1 next hop mask                 
    assign mgr_inst[47].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR47_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR47, Port2 next hop mask                 
    assign mgr_inst[47].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR47_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR47, Port3 next hop mask                 
    assign mgr_inst[47].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR47_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR48, Port0 next hop mask                 
    assign mgr_inst[48].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR48_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR48, Port1 next hop mask                 
    assign mgr_inst[48].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR48_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR48, Port2 next hop mask                 
    assign mgr_inst[48].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR48_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR48, Port3 next hop mask                 
    assign mgr_inst[48].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR48_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR49, Port0 next hop mask                 
    assign mgr_inst[49].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR49_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR49, Port1 next hop mask                 
    assign mgr_inst[49].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR49_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR49, Port2 next hop mask                 
    assign mgr_inst[49].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR49_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR49, Port3 next hop mask                 
    assign mgr_inst[49].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR49_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR50, Port0 next hop mask                 
    assign mgr_inst[50].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR50_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR50, Port1 next hop mask                 
    assign mgr_inst[50].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR50_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR50, Port2 next hop mask                 
    assign mgr_inst[50].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR50_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR50, Port3 next hop mask                 
    assign mgr_inst[50].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR50_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR51, Port0 next hop mask                 
    assign mgr_inst[51].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR51_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR51, Port1 next hop mask                 
    assign mgr_inst[51].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR51_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR51, Port2 next hop mask                 
    assign mgr_inst[51].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR51_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR51, Port3 next hop mask                 
    assign mgr_inst[51].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR51_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR52, Port0 next hop mask                 
    assign mgr_inst[52].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR52_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR52, Port1 next hop mask                 
    assign mgr_inst[52].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR52_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR52, Port2 next hop mask                 
    assign mgr_inst[52].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR52_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR52, Port3 next hop mask                 
    assign mgr_inst[52].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR52_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR53, Port0 next hop mask                 
    assign mgr_inst[53].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR53_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR53, Port1 next hop mask                 
    assign mgr_inst[53].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR53_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR53, Port2 next hop mask                 
    assign mgr_inst[53].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR53_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR53, Port3 next hop mask                 
    assign mgr_inst[53].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR53_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR54, Port0 next hop mask                 
    assign mgr_inst[54].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR54_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR54, Port1 next hop mask                 
    assign mgr_inst[54].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR54_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR54, Port2 next hop mask                 
    assign mgr_inst[54].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR54_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR54, Port3 next hop mask                 
    assign mgr_inst[54].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR54_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR55, Port0 next hop mask                 
    assign mgr_inst[55].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR55_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR55, Port1 next hop mask                 
    assign mgr_inst[55].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR55_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR55, Port2 next hop mask                 
    assign mgr_inst[55].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR55_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR55, Port3 next hop mask                 
    assign mgr_inst[55].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR55_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR56, Port0 next hop mask                 
    assign mgr_inst[56].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR56_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR56, Port1 next hop mask                 
    assign mgr_inst[56].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR56_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR56, Port2 next hop mask                 
    assign mgr_inst[56].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR56_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR56, Port3 next hop mask                 
    assign mgr_inst[56].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR56_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR57, Port0 next hop mask                 
    assign mgr_inst[57].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR57_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR57, Port1 next hop mask                 
    assign mgr_inst[57].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR57_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR57, Port2 next hop mask                 
    assign mgr_inst[57].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR57_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR57, Port3 next hop mask                 
    assign mgr_inst[57].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR57_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR58, Port0 next hop mask                 
    assign mgr_inst[58].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR58_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR58, Port1 next hop mask                 
    assign mgr_inst[58].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR58_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR58, Port2 next hop mask                 
    assign mgr_inst[58].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR58_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR58, Port3 next hop mask                 
    assign mgr_inst[58].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR58_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR59, Port0 next hop mask                 
    assign mgr_inst[59].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR59_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR59, Port1 next hop mask                 
    assign mgr_inst[59].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR59_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR59, Port2 next hop mask                 
    assign mgr_inst[59].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR59_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR59, Port3 next hop mask                 
    assign mgr_inst[59].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR59_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR60, Port0 next hop mask                 
    assign mgr_inst[60].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR60_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR60, Port1 next hop mask                 
    assign mgr_inst[60].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR60_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR60, Port2 next hop mask                 
    assign mgr_inst[60].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR60_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR60, Port3 next hop mask                 
    assign mgr_inst[60].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR60_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR61, Port0 next hop mask                 
    assign mgr_inst[61].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR61_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR61, Port1 next hop mask                 
    assign mgr_inst[61].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR61_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR61, Port2 next hop mask                 
    assign mgr_inst[61].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR61_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR61, Port3 next hop mask                 
    assign mgr_inst[61].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR61_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR62, Port0 next hop mask                 
    assign mgr_inst[62].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR62_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR62, Port1 next hop mask                 
    assign mgr_inst[62].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR62_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR62, Port2 next hop mask                 
    assign mgr_inst[62].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR62_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR62, Port3 next hop mask                 
    assign mgr_inst[62].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR62_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR63, Port0 next hop mask                 
    assign mgr_inst[63].sys__mgr__port0_destinationMask    = `NOC_CONT_MGR63_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR63, Port1 next hop mask                 
    assign mgr_inst[63].sys__mgr__port1_destinationMask    = `NOC_CONT_MGR63_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR63, Port2 next hop mask                 
    assign mgr_inst[63].sys__mgr__port2_destinationMask    = `NOC_CONT_MGR63_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR63, Port3 next hop mask                 
    assign mgr_inst[63].sys__mgr__port3_destinationMask    = `NOC_CONT_MGR63_PORT3_DESTINATION_MGR_BITMASK ;