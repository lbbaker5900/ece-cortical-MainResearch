
          assign read_ready_strm0   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM0_READ_ACCESS)  ;
          assign write_ready_strm0  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM0_WRITE_ACCESS) ;
          assign read_ready_strm1   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM1_READ_ACCESS)  ;
          assign write_ready_strm1  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM1_WRITE_ACCESS) ;
          assign read_ready_strm2   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM2_READ_ACCESS)  ;
          assign write_ready_strm2  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM2_WRITE_ACCESS) ;
          assign read_ready_strm3   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM3_READ_ACCESS)  ;
          assign write_ready_strm3  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM3_WRITE_ACCESS) ;
          assign read_ready_strm4   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM4_READ_ACCESS)  ;
          assign write_ready_strm4  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM4_WRITE_ACCESS) ;
          assign read_ready_strm5   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM5_READ_ACCESS)  ;
          assign write_ready_strm5  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM5_WRITE_ACCESS) ;
          assign read_ready_strm6   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM6_READ_ACCESS)  ;
          assign write_ready_strm6  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM6_WRITE_ACCESS) ;
          assign read_ready_strm7   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM7_READ_ACCESS)  ;
          assign write_ready_strm7  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM7_WRITE_ACCESS) ;
          assign read_ready_strm8   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM8_READ_ACCESS)  ;
          assign write_ready_strm8  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM8_WRITE_ACCESS) ;
          assign read_ready_strm9   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM9_READ_ACCESS)  ;
          assign write_ready_strm9  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM9_WRITE_ACCESS) ;
          assign read_ready_strm10   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM10_READ_ACCESS)  ;
          assign write_ready_strm10  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM10_WRITE_ACCESS) ;
          assign read_ready_strm11   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM11_READ_ACCESS)  ;
          assign write_ready_strm11  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM11_WRITE_ACCESS) ;
          assign read_ready_strm12   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM12_READ_ACCESS)  ;
          assign write_ready_strm12  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM12_WRITE_ACCESS) ;
          assign read_ready_strm13   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM13_READ_ACCESS)  ;
          assign write_ready_strm13  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM13_WRITE_ACCESS) ;
          assign read_ready_strm14   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM14_READ_ACCESS)  ;
          assign write_ready_strm14  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM14_WRITE_ACCESS) ;
          assign read_ready_strm15   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM15_READ_ACCESS)  ;
          assign write_ready_strm15  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM15_WRITE_ACCESS) ;
          assign read_ready_strm16   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM16_READ_ACCESS)  ;
          assign write_ready_strm16  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM16_WRITE_ACCESS) ;
          assign read_ready_strm17   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM17_READ_ACCESS)  ;
          assign write_ready_strm17  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM17_WRITE_ACCESS) ;
          assign read_ready_strm18   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM18_READ_ACCESS)  ;
          assign write_ready_strm18  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM18_WRITE_ACCESS) ;
          assign read_ready_strm19   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM19_READ_ACCESS)  ;
          assign write_ready_strm19  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM19_WRITE_ACCESS) ;
          assign read_ready_strm20   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM20_READ_ACCESS)  ;
          assign write_ready_strm20  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM20_WRITE_ACCESS) ;
          assign read_ready_strm21   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM21_READ_ACCESS)  ;
          assign write_ready_strm21  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM21_WRITE_ACCESS) ;
          assign read_ready_strm22   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM22_READ_ACCESS)  ;
          assign write_ready_strm22  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM22_WRITE_ACCESS) ;
          assign read_ready_strm23   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM23_READ_ACCESS)  ;
          assign write_ready_strm23  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM23_WRITE_ACCESS) ;
          assign read_ready_strm24   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM24_READ_ACCESS)  ;
          assign write_ready_strm24  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM24_WRITE_ACCESS) ;
          assign read_ready_strm25   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM25_READ_ACCESS)  ;
          assign write_ready_strm25  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM25_WRITE_ACCESS) ;
          assign read_ready_strm26   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM26_READ_ACCESS)  ;
          assign write_ready_strm26  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM26_WRITE_ACCESS) ;
          assign read_ready_strm27   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM27_READ_ACCESS)  ;
          assign write_ready_strm27  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM27_WRITE_ACCESS) ;
          assign read_ready_strm28   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM28_READ_ACCESS)  ;
          assign write_ready_strm28  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM28_WRITE_ACCESS) ;
          assign read_ready_strm29   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM29_READ_ACCESS)  ;
          assign write_ready_strm29  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM29_WRITE_ACCESS) ;
          assign read_ready_strm30   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM30_READ_ACCESS)  ;
          assign write_ready_strm30  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM30_WRITE_ACCESS) ;
          assign read_ready_strm31   = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM31_READ_ACCESS)  ;
          assign write_ready_strm31  = ( mem_acc_state_next == `MEM_ACC_CONT_DMA_STRM31_WRITE_ACCESS) ;