
  // NoC port 0
  output                                         mgr__noc__port0_valid           ;
  output   [`COMMON_STD_INTF_CNTL_RANGE       ]  mgr__noc__port0_cntl            ;
  output   [`MGR_NOC_CONT_NOC_PORT_DATA_RANGE ]  mgr__noc__port0_data            ;
  input                                          noc__mgr__port0_fc              ;
  input                                          noc__mgr__port0_valid           ;
  input    [`COMMON_STD_INTF_CNTL_RANGE       ]  noc__mgr__port0_cntl            ;
  input    [`MGR_NOC_CONT_NOC_PORT_DATA_RANGE ]  noc__mgr__port0_data            ;
  output                                         mgr__noc__port0_fc              ;
  input    [`MGR_HOST_MGR_ID_BITMASK_RANGE         ]  sys__mgr__port0_destinationMask ;

  // NoC port 1
  output                                         mgr__noc__port1_valid           ;
  output   [`COMMON_STD_INTF_CNTL_RANGE       ]  mgr__noc__port1_cntl            ;
  output   [`MGR_NOC_CONT_NOC_PORT_DATA_RANGE ]  mgr__noc__port1_data            ;
  input                                          noc__mgr__port1_fc              ;
  input                                          noc__mgr__port1_valid           ;
  input    [`COMMON_STD_INTF_CNTL_RANGE       ]  noc__mgr__port1_cntl            ;
  input    [`MGR_NOC_CONT_NOC_PORT_DATA_RANGE ]  noc__mgr__port1_data            ;
  output                                         mgr__noc__port1_fc              ;
  input    [`MGR_HOST_MGR_ID_BITMASK_RANGE         ]  sys__mgr__port1_destinationMask ;

  // NoC port 2
  output                                         mgr__noc__port2_valid           ;
  output   [`COMMON_STD_INTF_CNTL_RANGE       ]  mgr__noc__port2_cntl            ;
  output   [`MGR_NOC_CONT_NOC_PORT_DATA_RANGE ]  mgr__noc__port2_data            ;
  input                                          noc__mgr__port2_fc              ;
  input                                          noc__mgr__port2_valid           ;
  input    [`COMMON_STD_INTF_CNTL_RANGE       ]  noc__mgr__port2_cntl            ;
  input    [`MGR_NOC_CONT_NOC_PORT_DATA_RANGE ]  noc__mgr__port2_data            ;
  output                                         mgr__noc__port2_fc              ;
  input    [`MGR_HOST_MGR_ID_BITMASK_RANGE         ]  sys__mgr__port2_destinationMask ;

  // NoC port 3
  output                                         mgr__noc__port3_valid           ;
  output   [`COMMON_STD_INTF_CNTL_RANGE       ]  mgr__noc__port3_cntl            ;
  output   [`MGR_NOC_CONT_NOC_PORT_DATA_RANGE ]  mgr__noc__port3_data            ;
  input                                          noc__mgr__port3_fc              ;
  input                                          noc__mgr__port3_valid           ;
  input    [`COMMON_STD_INTF_CNTL_RANGE       ]  noc__mgr__port3_cntl            ;
  input    [`MGR_NOC_CONT_NOC_PORT_DATA_RANGE ]  noc__mgr__port3_data            ;
  output                                         mgr__noc__port3_fc              ;
  input    [`MGR_HOST_MGR_ID_BITMASK_RANGE         ]  sys__mgr__port3_destinationMask ;

