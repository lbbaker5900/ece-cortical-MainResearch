
  assign   mgr_inst[0].stu__mgr__valid     =   stu__mgr0__valid               ;
  assign   mgr_inst[0].stu__mgr__cntl      =   stu__mgr0__cntl                ;
  assign   mgr0__stu__ready                =   mgr_inst[0].mgr__stu__ready    ;
  assign   mgr_inst[0].stu__mgr__type      =   stu__mgr0__type                ;
  assign   mgr_inst[0].stu__mgr__data      =   stu__mgr0__data                ;
  assign   mgr_inst[0].stu__mgr__oob_data  =   stu__mgr0__oob_data            ;

  assign   mgr_inst[1].stu__mgr__valid     =   stu__mgr1__valid               ;
  assign   mgr_inst[1].stu__mgr__cntl      =   stu__mgr1__cntl                ;
  assign   mgr1__stu__ready                =   mgr_inst[1].mgr__stu__ready    ;
  assign   mgr_inst[1].stu__mgr__type      =   stu__mgr1__type                ;
  assign   mgr_inst[1].stu__mgr__data      =   stu__mgr1__data                ;
  assign   mgr_inst[1].stu__mgr__oob_data  =   stu__mgr1__oob_data            ;

  assign   mgr_inst[2].stu__mgr__valid     =   stu__mgr2__valid               ;
  assign   mgr_inst[2].stu__mgr__cntl      =   stu__mgr2__cntl                ;
  assign   mgr2__stu__ready                =   mgr_inst[2].mgr__stu__ready    ;
  assign   mgr_inst[2].stu__mgr__type      =   stu__mgr2__type                ;
  assign   mgr_inst[2].stu__mgr__data      =   stu__mgr2__data                ;
  assign   mgr_inst[2].stu__mgr__oob_data  =   stu__mgr2__oob_data            ;

  assign   mgr_inst[3].stu__mgr__valid     =   stu__mgr3__valid               ;
  assign   mgr_inst[3].stu__mgr__cntl      =   stu__mgr3__cntl                ;
  assign   mgr3__stu__ready                =   mgr_inst[3].mgr__stu__ready    ;
  assign   mgr_inst[3].stu__mgr__type      =   stu__mgr3__type                ;
  assign   mgr_inst[3].stu__mgr__data      =   stu__mgr3__data                ;
  assign   mgr_inst[3].stu__mgr__oob_data  =   stu__mgr3__oob_data            ;

