
  // General control and status                                                   
  input                                         mgr0__sys__allSynchronized     ;
  output                                        sys__mgr0__thisSynchronized    ;
  output                                        sys__mgr0__ready               ;
  output                                        sys__mgr0__complete            ;

  output                                        sys__pe0__allSynchronized     ;
  input                                         pe0__sys__thisSynchronized    ;
  input                                         pe0__sys__ready               ;
  input                                         pe0__sys__complete            ;

  // General control and status                                                   
  input                                         mgr1__sys__allSynchronized     ;
  output                                        sys__mgr1__thisSynchronized    ;
  output                                        sys__mgr1__ready               ;
  output                                        sys__mgr1__complete            ;

  output                                        sys__pe1__allSynchronized     ;
  input                                         pe1__sys__thisSynchronized    ;
  input                                         pe1__sys__ready               ;
  input                                         pe1__sys__complete            ;

  // General control and status                                                   
  input                                         mgr2__sys__allSynchronized     ;
  output                                        sys__mgr2__thisSynchronized    ;
  output                                        sys__mgr2__ready               ;
  output                                        sys__mgr2__complete            ;

  output                                        sys__pe2__allSynchronized     ;
  input                                         pe2__sys__thisSynchronized    ;
  input                                         pe2__sys__ready               ;
  input                                         pe2__sys__complete            ;

  // General control and status                                                   
  input                                         mgr3__sys__allSynchronized     ;
  output                                        sys__mgr3__thisSynchronized    ;
  output                                        sys__mgr3__ready               ;
  output                                        sys__mgr3__complete            ;

  output                                        sys__pe3__allSynchronized     ;
  input                                         pe3__sys__thisSynchronized    ;
  input                                         pe3__sys__ready               ;
  input                                         pe3__sys__complete            ;
