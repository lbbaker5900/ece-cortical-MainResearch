
      // Aggregate Control-path (cp) to NoC 
      noc__scntl__cp_ready      , 
      scntl__noc__cp_cntl       , 
      scntl__noc__cp_type       , 
      scntl__noc__cp_data       , 
      scntl__noc__cp_laneId     , 
      scntl__noc__cp_strmId     , 
      scntl__noc__cp_valid      , 
      // Aggregate Datapath (cp) from NoC 
      scntl__noc__cp_ready      , 
      noc__scntl__cp_cntl       , 
      noc__scntl__cp_type       , 
      noc__scntl__cp_data       , 
      noc__scntl__cp_peId       , 
      noc__scntl__cp_laneId     , 
      noc__scntl__cp_strmId     , 
      noc__scntl__cp_valid      , 

      // Aggregate Datapath (dp) to NoC 
      noc__scntl__dp_ready      , 
      scntl__noc__dp_cntl       , 
      scntl__noc__dp_type       , 
      scntl__noc__dp_peId       , 
      scntl__noc__dp_laneId     , 
      scntl__noc__dp_strmId     , 
      scntl__noc__dp_data       , 
      scntl__noc__dp_valid      , 
      // Aggregate Datapath (dp) from NoC 
      scntl__noc__dp_ready      , 
      noc__scntl__dp_cntl       , 
      noc__scntl__dp_type       , 
      noc__scntl__dp_laneId     , 
      noc__scntl__dp_strmId     , 
      noc__scntl__dp_data       , 
      noc__scntl__dp_valid      , 

      // Only one lane from each DMA can feed NoC
      // lane0 from NoC 
      sdp__cntl__lane0_strm_ready      , 
      cntl__sdp__lane0_strm_cntl       , 
      cntl__sdp__lane0_strm_id         , 
      cntl__sdp__lane0_strm_data       , 
      cntl__sdp__lane0_strm_data_valid , 
      // lane0 to NoC 
      cntl__sdp__lane0_strm_ready      , 
      sdp__cntl__lane0_strm_cntl       , 
      sdp__cntl__lane0_strm_id         , 
      sdp__cntl__lane0_strm_data       , 
      sdp__cntl__lane0_strm_data_valid , 
      // lane1 from NoC 
      sdp__cntl__lane1_strm_ready      , 
      cntl__sdp__lane1_strm_cntl       , 
      cntl__sdp__lane1_strm_id         , 
      cntl__sdp__lane1_strm_data       , 
      cntl__sdp__lane1_strm_data_valid , 
      // lane1 to NoC 
      cntl__sdp__lane1_strm_ready      , 
      sdp__cntl__lane1_strm_cntl       , 
      sdp__cntl__lane1_strm_id         , 
      sdp__cntl__lane1_strm_data       , 
      sdp__cntl__lane1_strm_data_valid , 
      // lane2 from NoC 
      sdp__cntl__lane2_strm_ready      , 
      cntl__sdp__lane2_strm_cntl       , 
      cntl__sdp__lane2_strm_id         , 
      cntl__sdp__lane2_strm_data       , 
      cntl__sdp__lane2_strm_data_valid , 
      // lane2 to NoC 
      cntl__sdp__lane2_strm_ready      , 
      sdp__cntl__lane2_strm_cntl       , 
      sdp__cntl__lane2_strm_id         , 
      sdp__cntl__lane2_strm_data       , 
      sdp__cntl__lane2_strm_data_valid , 
      // lane3 from NoC 
      sdp__cntl__lane3_strm_ready      , 
      cntl__sdp__lane3_strm_cntl       , 
      cntl__sdp__lane3_strm_id         , 
      cntl__sdp__lane3_strm_data       , 
      cntl__sdp__lane3_strm_data_valid , 
      // lane3 to NoC 
      cntl__sdp__lane3_strm_ready      , 
      sdp__cntl__lane3_strm_cntl       , 
      sdp__cntl__lane3_strm_id         , 
      sdp__cntl__lane3_strm_data       , 
      sdp__cntl__lane3_strm_data_valid , 
      // lane4 from NoC 
      sdp__cntl__lane4_strm_ready      , 
      cntl__sdp__lane4_strm_cntl       , 
      cntl__sdp__lane4_strm_id         , 
      cntl__sdp__lane4_strm_data       , 
      cntl__sdp__lane4_strm_data_valid , 
      // lane4 to NoC 
      cntl__sdp__lane4_strm_ready      , 
      sdp__cntl__lane4_strm_cntl       , 
      sdp__cntl__lane4_strm_id         , 
      sdp__cntl__lane4_strm_data       , 
      sdp__cntl__lane4_strm_data_valid , 
      // lane5 from NoC 
      sdp__cntl__lane5_strm_ready      , 
      cntl__sdp__lane5_strm_cntl       , 
      cntl__sdp__lane5_strm_id         , 
      cntl__sdp__lane5_strm_data       , 
      cntl__sdp__lane5_strm_data_valid , 
      // lane5 to NoC 
      cntl__sdp__lane5_strm_ready      , 
      sdp__cntl__lane5_strm_cntl       , 
      sdp__cntl__lane5_strm_id         , 
      sdp__cntl__lane5_strm_data       , 
      sdp__cntl__lane5_strm_data_valid , 
      // lane6 from NoC 
      sdp__cntl__lane6_strm_ready      , 
      cntl__sdp__lane6_strm_cntl       , 
      cntl__sdp__lane6_strm_id         , 
      cntl__sdp__lane6_strm_data       , 
      cntl__sdp__lane6_strm_data_valid , 
      // lane6 to NoC 
      cntl__sdp__lane6_strm_ready      , 
      sdp__cntl__lane6_strm_cntl       , 
      sdp__cntl__lane6_strm_id         , 
      sdp__cntl__lane6_strm_data       , 
      sdp__cntl__lane6_strm_data_valid , 
      // lane7 from NoC 
      sdp__cntl__lane7_strm_ready      , 
      cntl__sdp__lane7_strm_cntl       , 
      cntl__sdp__lane7_strm_id         , 
      cntl__sdp__lane7_strm_data       , 
      cntl__sdp__lane7_strm_data_valid , 
      // lane7 to NoC 
      cntl__sdp__lane7_strm_ready      , 
      sdp__cntl__lane7_strm_cntl       , 
      sdp__cntl__lane7_strm_id         , 
      sdp__cntl__lane7_strm_data       , 
      sdp__cntl__lane7_strm_data_valid , 
      // lane8 from NoC 
      sdp__cntl__lane8_strm_ready      , 
      cntl__sdp__lane8_strm_cntl       , 
      cntl__sdp__lane8_strm_id         , 
      cntl__sdp__lane8_strm_data       , 
      cntl__sdp__lane8_strm_data_valid , 
      // lane8 to NoC 
      cntl__sdp__lane8_strm_ready      , 
      sdp__cntl__lane8_strm_cntl       , 
      sdp__cntl__lane8_strm_id         , 
      sdp__cntl__lane8_strm_data       , 
      sdp__cntl__lane8_strm_data_valid , 
      // lane9 from NoC 
      sdp__cntl__lane9_strm_ready      , 
      cntl__sdp__lane9_strm_cntl       , 
      cntl__sdp__lane9_strm_id         , 
      cntl__sdp__lane9_strm_data       , 
      cntl__sdp__lane9_strm_data_valid , 
      // lane9 to NoC 
      cntl__sdp__lane9_strm_ready      , 
      sdp__cntl__lane9_strm_cntl       , 
      sdp__cntl__lane9_strm_id         , 
      sdp__cntl__lane9_strm_data       , 
      sdp__cntl__lane9_strm_data_valid , 
      // lane10 from NoC 
      sdp__cntl__lane10_strm_ready      , 
      cntl__sdp__lane10_strm_cntl       , 
      cntl__sdp__lane10_strm_id         , 
      cntl__sdp__lane10_strm_data       , 
      cntl__sdp__lane10_strm_data_valid , 
      // lane10 to NoC 
      cntl__sdp__lane10_strm_ready      , 
      sdp__cntl__lane10_strm_cntl       , 
      sdp__cntl__lane10_strm_id         , 
      sdp__cntl__lane10_strm_data       , 
      sdp__cntl__lane10_strm_data_valid , 
      // lane11 from NoC 
      sdp__cntl__lane11_strm_ready      , 
      cntl__sdp__lane11_strm_cntl       , 
      cntl__sdp__lane11_strm_id         , 
      cntl__sdp__lane11_strm_data       , 
      cntl__sdp__lane11_strm_data_valid , 
      // lane11 to NoC 
      cntl__sdp__lane11_strm_ready      , 
      sdp__cntl__lane11_strm_cntl       , 
      sdp__cntl__lane11_strm_id         , 
      sdp__cntl__lane11_strm_data       , 
      sdp__cntl__lane11_strm_data_valid , 
      // lane12 from NoC 
      sdp__cntl__lane12_strm_ready      , 
      cntl__sdp__lane12_strm_cntl       , 
      cntl__sdp__lane12_strm_id         , 
      cntl__sdp__lane12_strm_data       , 
      cntl__sdp__lane12_strm_data_valid , 
      // lane12 to NoC 
      cntl__sdp__lane12_strm_ready      , 
      sdp__cntl__lane12_strm_cntl       , 
      sdp__cntl__lane12_strm_id         , 
      sdp__cntl__lane12_strm_data       , 
      sdp__cntl__lane12_strm_data_valid , 
      // lane13 from NoC 
      sdp__cntl__lane13_strm_ready      , 
      cntl__sdp__lane13_strm_cntl       , 
      cntl__sdp__lane13_strm_id         , 
      cntl__sdp__lane13_strm_data       , 
      cntl__sdp__lane13_strm_data_valid , 
      // lane13 to NoC 
      cntl__sdp__lane13_strm_ready      , 
      sdp__cntl__lane13_strm_cntl       , 
      sdp__cntl__lane13_strm_id         , 
      sdp__cntl__lane13_strm_data       , 
      sdp__cntl__lane13_strm_data_valid , 
      // lane14 from NoC 
      sdp__cntl__lane14_strm_ready      , 
      cntl__sdp__lane14_strm_cntl       , 
      cntl__sdp__lane14_strm_id         , 
      cntl__sdp__lane14_strm_data       , 
      cntl__sdp__lane14_strm_data_valid , 
      // lane14 to NoC 
      cntl__sdp__lane14_strm_ready      , 
      sdp__cntl__lane14_strm_cntl       , 
      sdp__cntl__lane14_strm_id         , 
      sdp__cntl__lane14_strm_data       , 
      sdp__cntl__lane14_strm_data_valid , 
      // lane15 from NoC 
      sdp__cntl__lane15_strm_ready      , 
      cntl__sdp__lane15_strm_cntl       , 
      cntl__sdp__lane15_strm_id         , 
      cntl__sdp__lane15_strm_data       , 
      cntl__sdp__lane15_strm_data_valid , 
      // lane15 to NoC 
      cntl__sdp__lane15_strm_ready      , 
      sdp__cntl__lane15_strm_cntl       , 
      sdp__cntl__lane15_strm_id         , 
      sdp__cntl__lane15_strm_data       , 
      sdp__cntl__lane15_strm_data_valid , 
      // lane16 from NoC 
      sdp__cntl__lane16_strm_ready      , 
      cntl__sdp__lane16_strm_cntl       , 
      cntl__sdp__lane16_strm_id         , 
      cntl__sdp__lane16_strm_data       , 
      cntl__sdp__lane16_strm_data_valid , 
      // lane16 to NoC 
      cntl__sdp__lane16_strm_ready      , 
      sdp__cntl__lane16_strm_cntl       , 
      sdp__cntl__lane16_strm_id         , 
      sdp__cntl__lane16_strm_data       , 
      sdp__cntl__lane16_strm_data_valid , 
      // lane17 from NoC 
      sdp__cntl__lane17_strm_ready      , 
      cntl__sdp__lane17_strm_cntl       , 
      cntl__sdp__lane17_strm_id         , 
      cntl__sdp__lane17_strm_data       , 
      cntl__sdp__lane17_strm_data_valid , 
      // lane17 to NoC 
      cntl__sdp__lane17_strm_ready      , 
      sdp__cntl__lane17_strm_cntl       , 
      sdp__cntl__lane17_strm_id         , 
      sdp__cntl__lane17_strm_data       , 
      sdp__cntl__lane17_strm_data_valid , 
      // lane18 from NoC 
      sdp__cntl__lane18_strm_ready      , 
      cntl__sdp__lane18_strm_cntl       , 
      cntl__sdp__lane18_strm_id         , 
      cntl__sdp__lane18_strm_data       , 
      cntl__sdp__lane18_strm_data_valid , 
      // lane18 to NoC 
      cntl__sdp__lane18_strm_ready      , 
      sdp__cntl__lane18_strm_cntl       , 
      sdp__cntl__lane18_strm_id         , 
      sdp__cntl__lane18_strm_data       , 
      sdp__cntl__lane18_strm_data_valid , 
      // lane19 from NoC 
      sdp__cntl__lane19_strm_ready      , 
      cntl__sdp__lane19_strm_cntl       , 
      cntl__sdp__lane19_strm_id         , 
      cntl__sdp__lane19_strm_data       , 
      cntl__sdp__lane19_strm_data_valid , 
      // lane19 to NoC 
      cntl__sdp__lane19_strm_ready      , 
      sdp__cntl__lane19_strm_cntl       , 
      sdp__cntl__lane19_strm_id         , 
      sdp__cntl__lane19_strm_data       , 
      sdp__cntl__lane19_strm_data_valid , 
      // lane20 from NoC 
      sdp__cntl__lane20_strm_ready      , 
      cntl__sdp__lane20_strm_cntl       , 
      cntl__sdp__lane20_strm_id         , 
      cntl__sdp__lane20_strm_data       , 
      cntl__sdp__lane20_strm_data_valid , 
      // lane20 to NoC 
      cntl__sdp__lane20_strm_ready      , 
      sdp__cntl__lane20_strm_cntl       , 
      sdp__cntl__lane20_strm_id         , 
      sdp__cntl__lane20_strm_data       , 
      sdp__cntl__lane20_strm_data_valid , 
      // lane21 from NoC 
      sdp__cntl__lane21_strm_ready      , 
      cntl__sdp__lane21_strm_cntl       , 
      cntl__sdp__lane21_strm_id         , 
      cntl__sdp__lane21_strm_data       , 
      cntl__sdp__lane21_strm_data_valid , 
      // lane21 to NoC 
      cntl__sdp__lane21_strm_ready      , 
      sdp__cntl__lane21_strm_cntl       , 
      sdp__cntl__lane21_strm_id         , 
      sdp__cntl__lane21_strm_data       , 
      sdp__cntl__lane21_strm_data_valid , 
      // lane22 from NoC 
      sdp__cntl__lane22_strm_ready      , 
      cntl__sdp__lane22_strm_cntl       , 
      cntl__sdp__lane22_strm_id         , 
      cntl__sdp__lane22_strm_data       , 
      cntl__sdp__lane22_strm_data_valid , 
      // lane22 to NoC 
      cntl__sdp__lane22_strm_ready      , 
      sdp__cntl__lane22_strm_cntl       , 
      sdp__cntl__lane22_strm_id         , 
      sdp__cntl__lane22_strm_data       , 
      sdp__cntl__lane22_strm_data_valid , 
      // lane23 from NoC 
      sdp__cntl__lane23_strm_ready      , 
      cntl__sdp__lane23_strm_cntl       , 
      cntl__sdp__lane23_strm_id         , 
      cntl__sdp__lane23_strm_data       , 
      cntl__sdp__lane23_strm_data_valid , 
      // lane23 to NoC 
      cntl__sdp__lane23_strm_ready      , 
      sdp__cntl__lane23_strm_cntl       , 
      sdp__cntl__lane23_strm_id         , 
      sdp__cntl__lane23_strm_data       , 
      sdp__cntl__lane23_strm_data_valid , 
      // lane24 from NoC 
      sdp__cntl__lane24_strm_ready      , 
      cntl__sdp__lane24_strm_cntl       , 
      cntl__sdp__lane24_strm_id         , 
      cntl__sdp__lane24_strm_data       , 
      cntl__sdp__lane24_strm_data_valid , 
      // lane24 to NoC 
      cntl__sdp__lane24_strm_ready      , 
      sdp__cntl__lane24_strm_cntl       , 
      sdp__cntl__lane24_strm_id         , 
      sdp__cntl__lane24_strm_data       , 
      sdp__cntl__lane24_strm_data_valid , 
      // lane25 from NoC 
      sdp__cntl__lane25_strm_ready      , 
      cntl__sdp__lane25_strm_cntl       , 
      cntl__sdp__lane25_strm_id         , 
      cntl__sdp__lane25_strm_data       , 
      cntl__sdp__lane25_strm_data_valid , 
      // lane25 to NoC 
      cntl__sdp__lane25_strm_ready      , 
      sdp__cntl__lane25_strm_cntl       , 
      sdp__cntl__lane25_strm_id         , 
      sdp__cntl__lane25_strm_data       , 
      sdp__cntl__lane25_strm_data_valid , 
      // lane26 from NoC 
      sdp__cntl__lane26_strm_ready      , 
      cntl__sdp__lane26_strm_cntl       , 
      cntl__sdp__lane26_strm_id         , 
      cntl__sdp__lane26_strm_data       , 
      cntl__sdp__lane26_strm_data_valid , 
      // lane26 to NoC 
      cntl__sdp__lane26_strm_ready      , 
      sdp__cntl__lane26_strm_cntl       , 
      sdp__cntl__lane26_strm_id         , 
      sdp__cntl__lane26_strm_data       , 
      sdp__cntl__lane26_strm_data_valid , 
      // lane27 from NoC 
      sdp__cntl__lane27_strm_ready      , 
      cntl__sdp__lane27_strm_cntl       , 
      cntl__sdp__lane27_strm_id         , 
      cntl__sdp__lane27_strm_data       , 
      cntl__sdp__lane27_strm_data_valid , 
      // lane27 to NoC 
      cntl__sdp__lane27_strm_ready      , 
      sdp__cntl__lane27_strm_cntl       , 
      sdp__cntl__lane27_strm_id         , 
      sdp__cntl__lane27_strm_data       , 
      sdp__cntl__lane27_strm_data_valid , 
      // lane28 from NoC 
      sdp__cntl__lane28_strm_ready      , 
      cntl__sdp__lane28_strm_cntl       , 
      cntl__sdp__lane28_strm_id         , 
      cntl__sdp__lane28_strm_data       , 
      cntl__sdp__lane28_strm_data_valid , 
      // lane28 to NoC 
      cntl__sdp__lane28_strm_ready      , 
      sdp__cntl__lane28_strm_cntl       , 
      sdp__cntl__lane28_strm_id         , 
      sdp__cntl__lane28_strm_data       , 
      sdp__cntl__lane28_strm_data_valid , 
      // lane29 from NoC 
      sdp__cntl__lane29_strm_ready      , 
      cntl__sdp__lane29_strm_cntl       , 
      cntl__sdp__lane29_strm_id         , 
      cntl__sdp__lane29_strm_data       , 
      cntl__sdp__lane29_strm_data_valid , 
      // lane29 to NoC 
      cntl__sdp__lane29_strm_ready      , 
      sdp__cntl__lane29_strm_cntl       , 
      sdp__cntl__lane29_strm_id         , 
      sdp__cntl__lane29_strm_data       , 
      sdp__cntl__lane29_strm_data_valid , 
      // lane30 from NoC 
      sdp__cntl__lane30_strm_ready      , 
      cntl__sdp__lane30_strm_cntl       , 
      cntl__sdp__lane30_strm_id         , 
      cntl__sdp__lane30_strm_data       , 
      cntl__sdp__lane30_strm_data_valid , 
      // lane30 to NoC 
      cntl__sdp__lane30_strm_ready      , 
      sdp__cntl__lane30_strm_cntl       , 
      sdp__cntl__lane30_strm_id         , 
      sdp__cntl__lane30_strm_data       , 
      sdp__cntl__lane30_strm_data_valid , 
      // lane31 from NoC 
      sdp__cntl__lane31_strm_ready      , 
      cntl__sdp__lane31_strm_cntl       , 
      cntl__sdp__lane31_strm_id         , 
      cntl__sdp__lane31_strm_data       , 
      cntl__sdp__lane31_strm_data_valid , 
      // lane31 to NoC 
      cntl__sdp__lane31_strm_ready      , 
      sdp__cntl__lane31_strm_cntl       , 
      sdp__cntl__lane31_strm_id         , 
      sdp__cntl__lane31_strm_data       , 
      sdp__cntl__lane31_strm_data_valid , 
