
            .stu__mgr0__valid        ( stu__mgr0__valid     ),
            .stu__mgr0__cntl         ( stu__mgr0__cntl      ),
            .mgr0__stu__ready        ( mgr0__stu__ready     ),
            .stu__mgr0__type         ( stu__mgr0__type      ),
            .stu__mgr0__data         ( stu__mgr0__data      ),
            .stu__mgr0__oob_data     ( stu__mgr0__oob_data  ),

            .stu__mgr1__valid        ( stu__mgr1__valid     ),
            .stu__mgr1__cntl         ( stu__mgr1__cntl      ),
            .mgr1__stu__ready        ( mgr1__stu__ready     ),
            .stu__mgr1__type         ( stu__mgr1__type      ),
            .stu__mgr1__data         ( stu__mgr1__data      ),
            .stu__mgr1__oob_data     ( stu__mgr1__oob_data  ),

            .stu__mgr2__valid        ( stu__mgr2__valid     ),
            .stu__mgr2__cntl         ( stu__mgr2__cntl      ),
            .mgr2__stu__ready        ( mgr2__stu__ready     ),
            .stu__mgr2__type         ( stu__mgr2__type      ),
            .stu__mgr2__data         ( stu__mgr2__data      ),
            .stu__mgr2__oob_data     ( stu__mgr2__oob_data  ),

            .stu__mgr3__valid        ( stu__mgr3__valid     ),
            .stu__mgr3__cntl         ( stu__mgr3__cntl      ),
            .mgr3__stu__ready        ( mgr3__stu__ready     ),
            .stu__mgr3__type         ( stu__mgr3__type      ),
            .stu__mgr3__data         ( stu__mgr3__data      ),
            .stu__mgr3__oob_data     ( stu__mgr3__oob_data  ),

